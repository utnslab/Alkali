module __handler_OoO_DETECT_OoO_detection#()
(
	 input  wire clk, 
	 input  wire rst,
	//input ports STRUCT
	input wire [96-1:0] arg_28_tdata ,
	input wire  arg_28_tvalid ,
	output wire  arg_28_tready,
	//input ports BUF
	input wire [512-1:0] arg_29_tdata ,
	input wire [64-1:0] arg_29_tkeep ,
	input wire  arg_29_tlast ,
	input wire  arg_29_tvalid ,
	output wire  arg_29_tready,
	//input ports STRUCT
	input wire [184-1:0] arg_30_tdata ,
	input wire  arg_30_tvalid ,
	output wire  arg_30_tready,
	//input ports STRUCT
	input wire [112-1:0] arg_31_tdata ,
	input wire  arg_31_tvalid ,
	output wire  arg_31_tready,
	//input ports STRUCT
	input wire [160-1:0] arg_32_tdata ,
	input wire  arg_32_tvalid ,
	output wire  arg_32_tready,
	//output ports BUF
	output wire [512-1:0] DMA_WRITE_1_tdata ,
	output wire [64-1:0] DMA_WRITE_1_tkeep ,
	output wire  DMA_WRITE_1_tlast ,
	output wire  DMA_WRITE_1_tvalid ,
	input wire  DMA_WRITE_1_tready,
	//output ports STRUCT
	output wire [64-1:0] DMA_WRITE_2_tdata ,
	output wire  DMA_WRITE_2_tvalid ,
	input wire  DMA_WRITE_2_tready,
	//output ports BUF
	output wire [512-1:0] DMA_WRITE_3_tdata ,
	output wire [64-1:0] DMA_WRITE_3_tkeep ,
	output wire  DMA_WRITE_3_tlast ,
	output wire  DMA_WRITE_3_tvalid ,
	input wire  DMA_WRITE_3_tready,
	//output ports STRUCT
	output wire [184-1:0] DMA_WRITE_4_tdata ,
	output wire  DMA_WRITE_4_tvalid ,
	input wire  DMA_WRITE_4_tready,
	//output ports STRUCT
	output wire [112-1:0] DMA_WRITE_5_tdata ,
	output wire  DMA_WRITE_5_tvalid ,
	input wire  DMA_WRITE_5_tready,
	//output ports STRUCT
	output wire [160-1:0] DMA_WRITE_6_tdata ,
	output wire  DMA_WRITE_6_tvalid ,
	input wire  DMA_WRITE_6_tready,
	//output ports STRUCT
	output wire [96-1:0] outport_33_1_tdata ,
	output wire  outport_33_1_tvalid ,
	input wire  outport_33_1_tready,
	//output ports BUF
	output wire [512-1:0] outport_33_2_tdata ,
	output wire [64-1:0] outport_33_2_tkeep ,
	output wire  outport_33_2_tlast ,
	output wire  outport_33_2_tvalid ,
	input wire  outport_33_2_tready,
	//output ports STRUCT
	output wire [184-1:0] outport_33_3_tdata ,
	output wire  outport_33_3_tvalid ,
	input wire  outport_33_3_tready,
	//output ports STRUCT
	output wire [112-1:0] outport_33_4_tdata ,
	output wire  outport_33_4_tvalid ,
	input wire  outport_33_4_tready,
	//output ports STRUCT
	output wire [160-1:0] outport_33_5_tdata ,
	output wire  outport_33_5_tvalid ,
	input wire  outport_33_5_tready
);
//
 wire [96-1:0] arg_28_0_tdata;
 wire  arg_28_0_tvalid;
 wire  arg_28_0_tready;

//
 wire [96-1:0] arg_28_1_tdata;
 wire  arg_28_1_tvalid;
 wire  arg_28_1_tready;

//
 wire [96-1:0] arg_28_2_tdata;
 wire  arg_28_2_tvalid;
 wire  arg_28_2_tready;

axis_replication#(
.DATA_WIDTH(96),
.IF_STREAM(0),
.REAPLICA_COUNT(3)
)axis_replication_34(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.s_axis_in_tdata({arg_28_tdata}),
	.s_axis_in_tvalid({arg_28_tvalid}),
	.s_axis_in_tready({arg_28_tready}),
	//
	.m_axis_out_tdata({arg_28_0_tdata,arg_28_1_tdata,arg_28_2_tdata}),
	.m_axis_out_tvalid({arg_28_0_tvalid,arg_28_1_tvalid,arg_28_2_tvalid}),
	.m_axis_out_tready({arg_28_0_tready,arg_28_1_tready,arg_28_2_tready})
);

//
 wire [512-1:0] arg_29_0_tdata;
 wire [64-1:0] arg_29_0_tkeep;
 wire  arg_29_0_tvalid;
 wire  arg_29_0_tready;
 wire  arg_29_0_tlast;

//
 wire [512-1:0] arg_29_1_tdata;
 wire [64-1:0] arg_29_1_tkeep;
 wire  arg_29_1_tvalid;
 wire  arg_29_1_tready;
 wire  arg_29_1_tlast;

//
 wire [512-1:0] arg_29_2_tdata;
 wire [64-1:0] arg_29_2_tkeep;
 wire  arg_29_2_tvalid;
 wire  arg_29_2_tready;
 wire  arg_29_2_tlast;

axis_replication#(
.DATA_WIDTH(512),
.IF_STREAM(1),
.REAPLICA_COUNT(3)
)axis_replication_35(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.s_axis_in_tdata({arg_29_tdata}),
	.s_axis_in_tkeep({arg_29_tkeep}),
	.s_axis_in_tlast({arg_29_tlast}),
	.s_axis_in_tvalid({arg_29_tvalid}),
	.s_axis_in_tready({arg_29_tready}),
	//
	.m_axis_out_tdata({arg_29_0_tdata,arg_29_1_tdata,arg_29_2_tdata}),
	.m_axis_out_tkeep({arg_29_0_tkeep,arg_29_1_tkeep,arg_29_2_tkeep}),
	.m_axis_out_tlast({arg_29_0_tlast,arg_29_1_tlast,arg_29_2_tlast}),
	.m_axis_out_tvalid({arg_29_0_tvalid,arg_29_1_tvalid,arg_29_2_tvalid}),
	.m_axis_out_tready({arg_29_0_tready,arg_29_1_tready,arg_29_2_tready})
);

//
 wire [184-1:0] arg_30_0_tdata;
 wire  arg_30_0_tvalid;
 wire  arg_30_0_tready;

//
 wire [184-1:0] arg_30_1_tdata;
 wire  arg_30_1_tvalid;
 wire  arg_30_1_tready;

axis_replication#(
.DATA_WIDTH(184),
.IF_STREAM(0),
.REAPLICA_COUNT(2)
)axis_replication_36(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.s_axis_in_tdata({arg_30_tdata}),
	.s_axis_in_tvalid({arg_30_tvalid}),
	.s_axis_in_tready({arg_30_tready}),
	//
	.m_axis_out_tdata({arg_30_0_tdata,arg_30_1_tdata}),
	.m_axis_out_tvalid({arg_30_0_tvalid,arg_30_1_tvalid}),
	.m_axis_out_tready({arg_30_0_tready,arg_30_1_tready})
);

//
 wire [112-1:0] arg_31_0_tdata;
 wire  arg_31_0_tvalid;
 wire  arg_31_0_tready;

//
 wire [112-1:0] arg_31_1_tdata;
 wire  arg_31_1_tvalid;
 wire  arg_31_1_tready;

axis_replication#(
.DATA_WIDTH(112),
.IF_STREAM(0),
.REAPLICA_COUNT(2)
)axis_replication_37(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.s_axis_in_tdata({arg_31_tdata}),
	.s_axis_in_tvalid({arg_31_tvalid}),
	.s_axis_in_tready({arg_31_tready}),
	//
	.m_axis_out_tdata({arg_31_0_tdata,arg_31_1_tdata}),
	.m_axis_out_tvalid({arg_31_0_tvalid,arg_31_1_tvalid}),
	.m_axis_out_tready({arg_31_0_tready,arg_31_1_tready})
);

//
 wire [160-1:0] arg_32_0_tdata;
 wire  arg_32_0_tvalid;
 wire  arg_32_0_tready;

//
 wire [160-1:0] arg_32_1_tdata;
 wire  arg_32_1_tvalid;
 wire  arg_32_1_tready;

axis_replication#(
.DATA_WIDTH(160),
.IF_STREAM(0),
.REAPLICA_COUNT(2)
)axis_replication_38(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.s_axis_in_tdata({arg_32_tdata}),
	.s_axis_in_tvalid({arg_32_tvalid}),
	.s_axis_in_tready({arg_32_tready}),
	//
	.m_axis_out_tdata({arg_32_0_tdata,arg_32_1_tdata}),
	.m_axis_out_tvalid({arg_32_0_tvalid,arg_32_1_tvalid}),
	.m_axis_out_tready({arg_32_0_tready,arg_32_1_tready})
);

//const_INT
 wire [32-1:0] const_INT_39_tdata=0;
 wire  const_INT_39_tvalid=1;
 wire  const_INT_39_tready;

//const_INT
 wire [64-1:0] const_INT_40_tdata=0;
 wire  const_INT_40_tvalid=1;
 wire  const_INT_40_tready;

//Table lookup port wire def 
 wire [16-1:0] lookup_p_0_req_index;
 wire  lookup_p_0_req_valid;
 wire  lookup_p_0_req_ready;
 wire  lookup_p_0_value_valid;
 wire  lookup_p_0_value_ready;
 wire [256-1:0] lookup_p_0_value_data;

//Table update port wire def 
 wire [16-1:0] update_p_0_req_index;
 wire  update_p_0_req_index_valid;
 wire  update_p_0_req_index_ready;
 wire [256-1:0] update_p_0_req_data;
 wire  update_p_0_req_data_valid;
 wire  update_p_0_req_data_ready;

cam_arbiter#(
.TABLE_SIZE(16),
.KEY_SIZE(16),
.VALUE_SIZE(256),
.LOOKUP_PORTS(1),
.UPDATE_PORTS(1)
)table_41(
	 .clk(clk), 
	 .rst(rst) ,
	//lookup port 
	.s_lookup_req_index({lookup_p_0_req_index}),
	.s_lookup_req_valid({lookup_p_0_req_valid}),
	.s_lookup_req_ready({lookup_p_0_req_ready}),
	.s_lookup_value_valid({lookup_p_0_value_valid}),
	.s_lookup_value_data({lookup_p_0_value_data}),
	.s_lookup_value_ready({lookup_p_0_value_ready}),
	//update port 
	.s_update_req_index({update_p_0_req_index}),
	.s_update_req_index_valid({update_p_0_req_index_valid}),
	.s_update_req_index_ready({update_p_0_req_index_ready}),
	.s_update_req_data({update_p_0_req_data}),
	.s_update_req_data_valid({update_p_0_req_data_valid}),
	.s_update_req_data_ready({update_p_0_req_data_ready})
);

//Access Struct
 wire [32-1:0] struct_accessed_INT_43_tdata;
 wire  struct_accessed_INT_43_tvalid;
 wire  struct_accessed_INT_43_tready;

struct_access#(
.STRUCT_WIDTH(96),
.ACCESS_OFFSET(0),
.ACCESS_SIZE(32)
)struct_access_42(
	 .clk(clk), 
	 .rst(rst) ,
	//struct input
	.s_struct_axis_tdata({arg_28_0_tdata}),
	.s_struct_axis_tvalid({arg_28_0_tvalid}),
	.s_struct_axis_tready({arg_28_0_tready}),
	//output val
	.m_val_axis_tdata({struct_accessed_INT_43_tdata}),
	.m_val_axis_tvalid({struct_accessed_INT_43_tvalid}),
	.m_val_axis_tready({struct_accessed_INT_43_tready})
);

//bitcast dst
 wire [16-1:0] bitcasted_44_tdata;
 wire  bitcasted_44_tvalid;
 wire  bitcasted_44_tready;

//bitcast dst
 wire [16-1:0] bitcasted_44_0_tdata;
 wire  bitcasted_44_0_tvalid;
 wire  bitcasted_44_0_tready;

//bitcast dst
 wire [16-1:0] bitcasted_44_1_tdata;
 wire  bitcasted_44_1_tvalid;
 wire  bitcasted_44_1_tready;

axis_replication#(
.DATA_WIDTH(16),
.IF_STREAM(0),
.REAPLICA_COUNT(2)
)axis_replication_45(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.s_axis_in_tdata({bitcasted_44_tdata}),
	.s_axis_in_tvalid({bitcasted_44_tvalid}),
	.s_axis_in_tready({bitcasted_44_tready}),
	//
	.m_axis_out_tdata({bitcasted_44_0_tdata,bitcasted_44_1_tdata}),
	.m_axis_out_tvalid({bitcasted_44_0_tvalid,bitcasted_44_1_tvalid}),
	.m_axis_out_tready({bitcasted_44_0_tready,bitcasted_44_1_tready})
);

 assign bitcasted_44_tdata = struct_accessed_INT_43_tdata;
 assign bitcasted_44_tvalid = struct_accessed_INT_43_tvalid;
 assign struct_accessed_INT_43_tready = bitcasted_44_tready;

 assign lookup_p_0_req_index = bitcasted_44_0_tdata;
 assign lookup_p_0_req_valid = bitcasted_44_0_tvalid;
 assign bitcasted_44_0_tready = lookup_p_0_req_ready;

//table lookup resultlookedup_STRUCT_46
 wire [256-1:0] lookedup_STRUCT_46_tdata;
 wire  lookedup_STRUCT_46_tvalid;
 wire  lookedup_STRUCT_46_tready;

//table lookup resultlookedup_STRUCT_46
 wire [256-1:0] lookedup_STRUCT_46_0_tdata;
 wire  lookedup_STRUCT_46_0_tvalid;
 wire  lookedup_STRUCT_46_0_tready;

//table lookup resultlookedup_STRUCT_46
 wire [256-1:0] lookedup_STRUCT_46_1_tdata;
 wire  lookedup_STRUCT_46_1_tvalid;
 wire  lookedup_STRUCT_46_1_tready;

//table lookup resultlookedup_STRUCT_46
 wire [256-1:0] lookedup_STRUCT_46_2_tdata;
 wire  lookedup_STRUCT_46_2_tvalid;
 wire  lookedup_STRUCT_46_2_tready;

//table lookup resultlookedup_STRUCT_46
 wire [256-1:0] lookedup_STRUCT_46_3_tdata;
 wire  lookedup_STRUCT_46_3_tvalid;
 wire  lookedup_STRUCT_46_3_tready;

//table lookup resultlookedup_STRUCT_46
 wire [256-1:0] lookedup_STRUCT_46_4_tdata;
 wire  lookedup_STRUCT_46_4_tvalid;
 wire  lookedup_STRUCT_46_4_tready;

axis_replication#(
.DATA_WIDTH(256),
.IF_STREAM(0),
.REAPLICA_COUNT(5)
)axis_replication_47(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.s_axis_in_tdata({lookedup_STRUCT_46_tdata}),
	.s_axis_in_tvalid({lookedup_STRUCT_46_tvalid}),
	.s_axis_in_tready({lookedup_STRUCT_46_tready}),
	//
	.m_axis_out_tdata({lookedup_STRUCT_46_0_tdata,lookedup_STRUCT_46_1_tdata,lookedup_STRUCT_46_2_tdata,lookedup_STRUCT_46_3_tdata,lookedup_STRUCT_46_4_tdata}),
	.m_axis_out_tvalid({lookedup_STRUCT_46_0_tvalid,lookedup_STRUCT_46_1_tvalid,lookedup_STRUCT_46_2_tvalid,lookedup_STRUCT_46_3_tvalid,lookedup_STRUCT_46_4_tvalid}),
	.m_axis_out_tready({lookedup_STRUCT_46_0_tready,lookedup_STRUCT_46_1_tready,lookedup_STRUCT_46_2_tready,lookedup_STRUCT_46_3_tready,lookedup_STRUCT_46_4_tready})
);

 assign lookedup_STRUCT_46_tdata = lookup_p_0_value_data;
 assign lookedup_STRUCT_46_tvalid = lookup_p_0_value_valid;
 assign lookup_p_0_value_ready = lookedup_STRUCT_46_tready;

//inited_STRUCT
 wire [64-1:0] inited_STRUCT_48_tdata=0;
 wire  inited_STRUCT_48_tvalid=1;
 wire  inited_STRUCT_48_tready;

//inited_STRUCT
 wire [96-1:0] inited_STRUCT_49_tdata=0;
 wire  inited_STRUCT_49_tvalid=1;
 wire  inited_STRUCT_49_tready;

//Access Struct
 wire [32-1:0] struct_accessed_INT_51_tdata;
 wire  struct_accessed_INT_51_tvalid;
 wire  struct_accessed_INT_51_tready;

struct_access#(
.STRUCT_WIDTH(256),
.ACCESS_OFFSET(128),
.ACCESS_SIZE(32)
)struct_access_50(
	 .clk(clk), 
	 .rst(rst) ,
	//struct input
	.s_struct_axis_tdata({lookedup_STRUCT_46_0_tdata}),
	.s_struct_axis_tvalid({lookedup_STRUCT_46_0_tvalid}),
	.s_struct_axis_tready({lookedup_STRUCT_46_0_tready}),
	//output val
	.m_val_axis_tdata({struct_accessed_INT_51_tdata}),
	.m_val_axis_tvalid({struct_accessed_INT_51_tvalid}),
	.m_val_axis_tready({struct_accessed_INT_51_tready})
);

//Access Struct
 wire [32-1:0] struct_accessed_INT_53_tdata;
 wire  struct_accessed_INT_53_tvalid;
 wire  struct_accessed_INT_53_tready;

struct_access#(
.STRUCT_WIDTH(96),
.ACCESS_OFFSET(64),
.ACCESS_SIZE(32)
)struct_access_52(
	 .clk(clk), 
	 .rst(rst) ,
	//struct input
	.s_struct_axis_tdata({arg_28_1_tdata}),
	.s_struct_axis_tvalid({arg_28_1_tvalid}),
	.s_struct_axis_tready({arg_28_1_tready}),
	//output val
	.m_val_axis_tdata({struct_accessed_INT_53_tdata}),
	.m_val_axis_tvalid({struct_accessed_INT_53_tvalid}),
	.m_val_axis_tready({struct_accessed_INT_53_tready})
);

//Arithmetic OP Out
 wire [32-1:0] SUB_54_out_INT_55_tdata;
 wire  SUB_54_out_INT_55_tvalid;
 wire  SUB_54_out_INT_55_tready;

//Arithmetic OP Out
 wire [32-1:0] SUB_54_out_INT_55_0_tdata;
 wire  SUB_54_out_INT_55_0_tvalid;
 wire  SUB_54_out_INT_55_0_tready;

//Arithmetic OP Out
 wire [32-1:0] SUB_54_out_INT_55_1_tdata;
 wire  SUB_54_out_INT_55_1_tvalid;
 wire  SUB_54_out_INT_55_1_tready;

//Arithmetic OP Out
 wire [32-1:0] SUB_54_out_INT_55_2_tdata;
 wire  SUB_54_out_INT_55_2_tvalid;
 wire  SUB_54_out_INT_55_2_tready;

axis_replication#(
.DATA_WIDTH(32),
.IF_STREAM(0),
.REAPLICA_COUNT(3)
)axis_replication_56(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.s_axis_in_tdata({SUB_54_out_INT_55_tdata}),
	.s_axis_in_tvalid({SUB_54_out_INT_55_tvalid}),
	.s_axis_in_tready({SUB_54_out_INT_55_tready}),
	//
	.m_axis_out_tdata({SUB_54_out_INT_55_0_tdata,SUB_54_out_INT_55_1_tdata,SUB_54_out_INT_55_2_tdata}),
	.m_axis_out_tvalid({SUB_54_out_INT_55_0_tvalid,SUB_54_out_INT_55_1_tvalid,SUB_54_out_INT_55_2_tvalid}),
	.m_axis_out_tready({SUB_54_out_INT_55_0_tready,SUB_54_out_INT_55_1_tready,SUB_54_out_INT_55_2_tready})
);

ALU#(
.LVAL_SIZE(32),
.RVAL_SIZE(32),
.RESULT_SIZE(32),
.OPID(0)
)SUB_54(
	 .clk(clk), 
	 .rst(rst) ,
	//lval input
	.s_lval_axis_tdata({struct_accessed_INT_51_tdata}),
	.s_lval_axis_tvalid({struct_accessed_INT_51_tvalid}),
	.s_lval_axis_tready({struct_accessed_INT_51_tready}),
	//rval input
	.s_rval_axis_tdata({struct_accessed_INT_53_tdata}),
	.s_rval_axis_tvalid({struct_accessed_INT_53_tvalid}),
	.s_rval_axis_tready({struct_accessed_INT_53_tready}),
	//output val
	.m_val_axis_tdata({SUB_54_out_INT_55_tdata}),
	.m_val_axis_tvalid({SUB_54_out_INT_55_tvalid}),
	.m_val_axis_tready({SUB_54_out_INT_55_tready})
);

//Access Struct
 wire [32-1:0] struct_accessed_INT_58_tdata;
 wire  struct_accessed_INT_58_tvalid;
 wire  struct_accessed_INT_58_tready;

//Access Struct
 wire [32-1:0] struct_accessed_INT_58_0_tdata;
 wire  struct_accessed_INT_58_0_tvalid;
 wire  struct_accessed_INT_58_0_tready;

//Access Struct
 wire [32-1:0] struct_accessed_INT_58_1_tdata;
 wire  struct_accessed_INT_58_1_tvalid;
 wire  struct_accessed_INT_58_1_tready;

//Access Struct
 wire [32-1:0] struct_accessed_INT_58_2_tdata;
 wire  struct_accessed_INT_58_2_tvalid;
 wire  struct_accessed_INT_58_2_tready;

axis_replication#(
.DATA_WIDTH(32),
.IF_STREAM(0),
.REAPLICA_COUNT(3)
)axis_replication_59(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.s_axis_in_tdata({struct_accessed_INT_58_tdata}),
	.s_axis_in_tvalid({struct_accessed_INT_58_tvalid}),
	.s_axis_in_tready({struct_accessed_INT_58_tready}),
	//
	.m_axis_out_tdata({struct_accessed_INT_58_0_tdata,struct_accessed_INT_58_1_tdata,struct_accessed_INT_58_2_tdata}),
	.m_axis_out_tvalid({struct_accessed_INT_58_0_tvalid,struct_accessed_INT_58_1_tvalid,struct_accessed_INT_58_2_tvalid}),
	.m_axis_out_tready({struct_accessed_INT_58_0_tready,struct_accessed_INT_58_1_tready,struct_accessed_INT_58_2_tready})
);

struct_access#(
.STRUCT_WIDTH(96),
.ACCESS_OFFSET(32),
.ACCESS_SIZE(32)
)struct_access_57(
	 .clk(clk), 
	 .rst(rst) ,
	//struct input
	.s_struct_axis_tdata({arg_28_2_tdata}),
	.s_struct_axis_tvalid({arg_28_2_tvalid}),
	.s_struct_axis_tready({arg_28_2_tready}),
	//output val
	.m_val_axis_tdata({struct_accessed_INT_58_tdata}),
	.m_val_axis_tvalid({struct_accessed_INT_58_tvalid}),
	.m_val_axis_tready({struct_accessed_INT_58_tready})
);

//Arithmetic OP Out
 wire [32-1:0] SUB_60_out_INT_61_tdata;
 wire  SUB_60_out_INT_61_tvalid;
 wire  SUB_60_out_INT_61_tready;

//Arithmetic OP Out
 wire [32-1:0] SUB_60_out_INT_61_0_tdata;
 wire  SUB_60_out_INT_61_0_tvalid;
 wire  SUB_60_out_INT_61_0_tready;

//Arithmetic OP Out
 wire [32-1:0] SUB_60_out_INT_61_1_tdata;
 wire  SUB_60_out_INT_61_1_tvalid;
 wire  SUB_60_out_INT_61_1_tready;

axis_replication#(
.DATA_WIDTH(32),
.IF_STREAM(0),
.REAPLICA_COUNT(2)
)axis_replication_62(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.s_axis_in_tdata({SUB_60_out_INT_61_tdata}),
	.s_axis_in_tvalid({SUB_60_out_INT_61_tvalid}),
	.s_axis_in_tready({SUB_60_out_INT_61_tready}),
	//
	.m_axis_out_tdata({SUB_60_out_INT_61_0_tdata,SUB_60_out_INT_61_1_tdata}),
	.m_axis_out_tvalid({SUB_60_out_INT_61_0_tvalid,SUB_60_out_INT_61_1_tvalid}),
	.m_axis_out_tready({SUB_60_out_INT_61_0_tready,SUB_60_out_INT_61_1_tready})
);

ALU#(
.LVAL_SIZE(32),
.RVAL_SIZE(32),
.RESULT_SIZE(32),
.OPID(0)
)SUB_60(
	 .clk(clk), 
	 .rst(rst) ,
	//lval input
	.s_lval_axis_tdata({struct_accessed_INT_58_0_tdata}),
	.s_lval_axis_tvalid({struct_accessed_INT_58_0_tvalid}),
	.s_lval_axis_tready({struct_accessed_INT_58_0_tready}),
	//rval input
	.s_rval_axis_tdata({SUB_54_out_INT_55_0_tdata}),
	.s_rval_axis_tvalid({SUB_54_out_INT_55_0_tvalid}),
	.s_rval_axis_tready({SUB_54_out_INT_55_0_tready}),
	//output val
	.m_val_axis_tdata({SUB_60_out_INT_61_tdata}),
	.m_val_axis_tvalid({SUB_60_out_INT_61_tvalid}),
	.m_val_axis_tready({SUB_60_out_INT_61_tready})
);

//Access Struct
 wire [32-1:0] struct_accessed_INT_64_tdata;
 wire  struct_accessed_INT_64_tvalid;
 wire  struct_accessed_INT_64_tready;

//Access Struct
 wire [32-1:0] struct_accessed_INT_64_0_tdata;
 wire  struct_accessed_INT_64_0_tvalid;
 wire  struct_accessed_INT_64_0_tready;

//Access Struct
 wire [32-1:0] struct_accessed_INT_64_1_tdata;
 wire  struct_accessed_INT_64_1_tvalid;
 wire  struct_accessed_INT_64_1_tready;

//Access Struct
 wire [32-1:0] struct_accessed_INT_64_2_tdata;
 wire  struct_accessed_INT_64_2_tvalid;
 wire  struct_accessed_INT_64_2_tready;

axis_replication#(
.DATA_WIDTH(32),
.IF_STREAM(0),
.REAPLICA_COUNT(3)
)axis_replication_65(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.s_axis_in_tdata({struct_accessed_INT_64_tdata}),
	.s_axis_in_tvalid({struct_accessed_INT_64_tvalid}),
	.s_axis_in_tready({struct_accessed_INT_64_tready}),
	//
	.m_axis_out_tdata({struct_accessed_INT_64_0_tdata,struct_accessed_INT_64_1_tdata,struct_accessed_INT_64_2_tdata}),
	.m_axis_out_tvalid({struct_accessed_INT_64_0_tvalid,struct_accessed_INT_64_1_tvalid,struct_accessed_INT_64_2_tvalid}),
	.m_axis_out_tready({struct_accessed_INT_64_0_tready,struct_accessed_INT_64_1_tready,struct_accessed_INT_64_2_tready})
);

struct_access#(
.STRUCT_WIDTH(256),
.ACCESS_OFFSET(96),
.ACCESS_SIZE(32)
)struct_access_63(
	 .clk(clk), 
	 .rst(rst) ,
	//struct input
	.s_struct_axis_tdata({lookedup_STRUCT_46_1_tdata}),
	.s_struct_axis_tvalid({lookedup_STRUCT_46_1_tvalid}),
	.s_struct_axis_tready({lookedup_STRUCT_46_1_tready}),
	//output val
	.m_val_axis_tdata({struct_accessed_INT_64_tdata}),
	.m_val_axis_tvalid({struct_accessed_INT_64_tvalid}),
	.m_val_axis_tready({struct_accessed_INT_64_tready})
);

//Arithmetic OP Out
 wire [1-1:0] LT_66_out_INT_67_tdata;
 wire  LT_66_out_INT_67_tvalid;
 wire  LT_66_out_INT_67_tready;

ALU#(
.LVAL_SIZE(32),
.RVAL_SIZE(32),
.RESULT_SIZE(1),
.OPID(3)
)LT_66(
	 .clk(clk), 
	 .rst(rst) ,
	//lval input
	.s_lval_axis_tdata({SUB_60_out_INT_61_0_tdata}),
	.s_lval_axis_tvalid({SUB_60_out_INT_61_0_tvalid}),
	.s_lval_axis_tready({SUB_60_out_INT_61_0_tready}),
	//rval input
	.s_rval_axis_tdata({struct_accessed_INT_64_0_tdata}),
	.s_rval_axis_tvalid({struct_accessed_INT_64_0_tvalid}),
	.s_rval_axis_tready({struct_accessed_INT_64_0_tready}),
	//output val
	.m_val_axis_tdata({LT_66_out_INT_67_tdata}),
	.m_val_axis_tvalid({LT_66_out_INT_67_tvalid}),
	.m_val_axis_tready({LT_66_out_INT_67_tready})
);

//Arithmetic OP Out
 wire [32-1:0] SUB_68_out_INT_69_tdata;
 wire  SUB_68_out_INT_69_tvalid;
 wire  SUB_68_out_INT_69_tready;

ALU#(
.LVAL_SIZE(32),
.RVAL_SIZE(32),
.RESULT_SIZE(32),
.OPID(0)
)SUB_68(
	 .clk(clk), 
	 .rst(rst) ,
	//lval input
	.s_lval_axis_tdata({SUB_60_out_INT_61_1_tdata}),
	.s_lval_axis_tvalid({SUB_60_out_INT_61_1_tvalid}),
	.s_lval_axis_tready({SUB_60_out_INT_61_1_tready}),
	//rval input
	.s_rval_axis_tdata({struct_accessed_INT_64_1_tdata}),
	.s_rval_axis_tvalid({struct_accessed_INT_64_1_tvalid}),
	.s_rval_axis_tready({struct_accessed_INT_64_1_tready}),
	//output val
	.m_val_axis_tdata({SUB_68_out_INT_69_tdata}),
	.m_val_axis_tvalid({SUB_68_out_INT_69_tvalid}),
	.m_val_axis_tready({SUB_68_out_INT_69_tready})
);

//Arithmetic OP Out
 wire [1-1:0] LE_70_out_INT_71_tdata;
 wire  LE_70_out_INT_71_tvalid;
 wire  LE_70_out_INT_71_tready;

//Arithmetic OP Out
 wire [1-1:0] LE_70_out_INT_71_0_tdata;
 wire  LE_70_out_INT_71_0_tvalid;
 wire  LE_70_out_INT_71_0_tready;

//Arithmetic OP Out
 wire [1-1:0] LE_70_out_INT_71_1_tdata;
 wire  LE_70_out_INT_71_1_tvalid;
 wire  LE_70_out_INT_71_1_tready;

//Arithmetic OP Out
 wire [1-1:0] LE_70_out_INT_71_2_tdata;
 wire  LE_70_out_INT_71_2_tvalid;
 wire  LE_70_out_INT_71_2_tready;

axis_replication#(
.DATA_WIDTH(1),
.IF_STREAM(0),
.REAPLICA_COUNT(3)
)axis_replication_72(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.s_axis_in_tdata({LE_70_out_INT_71_tdata}),
	.s_axis_in_tvalid({LE_70_out_INT_71_tvalid}),
	.s_axis_in_tready({LE_70_out_INT_71_tready}),
	//
	.m_axis_out_tdata({LE_70_out_INT_71_0_tdata,LE_70_out_INT_71_1_tdata,LE_70_out_INT_71_2_tdata}),
	.m_axis_out_tvalid({LE_70_out_INT_71_0_tvalid,LE_70_out_INT_71_1_tvalid,LE_70_out_INT_71_2_tvalid}),
	.m_axis_out_tready({LE_70_out_INT_71_0_tready,LE_70_out_INT_71_1_tready,LE_70_out_INT_71_2_tready})
);

ALU#(
.LVAL_SIZE(32),
.RVAL_SIZE(32),
.RESULT_SIZE(1),
.OPID(6)
)LE_70(
	 .clk(clk), 
	 .rst(rst) ,
	//lval input
	.s_lval_axis_tdata({SUB_54_out_INT_55_1_tdata}),
	.s_lval_axis_tvalid({SUB_54_out_INT_55_1_tvalid}),
	.s_lval_axis_tready({SUB_54_out_INT_55_1_tready}),
	//rval input
	.s_rval_axis_tdata({struct_accessed_INT_58_1_tdata}),
	.s_rval_axis_tvalid({struct_accessed_INT_58_1_tvalid}),
	.s_rval_axis_tready({struct_accessed_INT_58_1_tready}),
	//output val
	.m_val_axis_tdata({LE_70_out_INT_71_tdata}),
	.m_val_axis_tvalid({LE_70_out_INT_71_tvalid}),
	.m_val_axis_tready({LE_70_out_INT_71_tready})
);

//Access Struct
 wire [32-1:0] struct_accessed_INT_74_tdata;
 wire  struct_accessed_INT_74_tvalid;
 wire  struct_accessed_INT_74_tready;

struct_access#(
.STRUCT_WIDTH(256),
.ACCESS_OFFSET(160),
.ACCESS_SIZE(32)
)struct_access_73(
	 .clk(clk), 
	 .rst(rst) ,
	//struct input
	.s_struct_axis_tdata({lookedup_STRUCT_46_2_tdata}),
	.s_struct_axis_tvalid({lookedup_STRUCT_46_2_tvalid}),
	.s_struct_axis_tready({lookedup_STRUCT_46_2_tready}),
	//output val
	.m_val_axis_tdata({struct_accessed_INT_74_tdata}),
	.m_val_axis_tvalid({struct_accessed_INT_74_tvalid}),
	.m_val_axis_tready({struct_accessed_INT_74_tready})
);

//struct_assign_75 output struct
 wire [64-1:0] structvar_76_tdata;
 wire  structvar_76_tvalid;
 wire  structvar_76_tready;

struct_assign#(
.STRUCT_WIDTH(64),
.ASSIGN_OFFSET(0),
.ASSIGN_SIZE(32)
)struct_assign_75(
	 .clk(clk), 
	 .rst(rst) ,
	//input struct
	.s_struct_axis_tdata({inited_STRUCT_48_tdata}),
	.s_struct_axis_tvalid({inited_STRUCT_48_tvalid}),
	.s_struct_axis_tready({inited_STRUCT_48_tready}),
	//input val
	.s_assignv_axis_tdata({struct_accessed_INT_74_tdata}),
	.s_assignv_axis_tvalid({struct_accessed_INT_74_tvalid}),
	.s_assignv_axis_tready({struct_accessed_INT_74_tready}),
	//output struct
	.m_struct_axis_tdata({structvar_76_tdata}),
	.m_struct_axis_tvalid({structvar_76_tvalid}),
	.m_struct_axis_tready({structvar_76_tready})
);

//
 wire [32-1:0] select_result_77_tdata;
 wire  select_result_77_tvalid;
 wire  select_result_77_tready;

select#(
.VAL_WIDTH(32),
.COND_WIDTH(1)
)select_78(
	 .clk(clk), 
	 .rst(rst) ,
	//select condition
	.s_cond_axis_tdata({LT_66_out_INT_67_tdata}),
	.s_cond_axis_tvalid({LT_66_out_INT_67_tvalid}),
	.s_cond_axis_tready({LT_66_out_INT_67_tready}),
	//select true val
	.s_true_val_axis_tdata({const_INT_39_tdata}),
	.s_true_val_axis_tvalid({const_INT_39_tvalid}),
	.s_true_val_axis_tready({const_INT_39_tready}),
	//select false val
	.s_false_val_axis_tdata({SUB_68_out_INT_69_tdata}),
	.s_false_val_axis_tvalid({SUB_68_out_INT_69_tvalid}),
	.s_false_val_axis_tready({SUB_68_out_INT_69_tready}),
	//select result
	.m_val_axis_tdata({select_result_77_tdata}),
	.m_val_axis_tvalid({select_result_77_tvalid}),
	.m_val_axis_tready({select_result_77_tready})
);

//Arithmetic OP Out
 wire [32-1:0] ADD_79_out_INT_80_tdata;
 wire  ADD_79_out_INT_80_tvalid;
 wire  ADD_79_out_INT_80_tready;

ALU#(
.LVAL_SIZE(32),
.RVAL_SIZE(32),
.RESULT_SIZE(32),
.OPID(1)
)ADD_79(
	 .clk(clk), 
	 .rst(rst) ,
	//lval input
	.s_lval_axis_tdata({SUB_54_out_INT_55_2_tdata}),
	.s_lval_axis_tvalid({SUB_54_out_INT_55_2_tvalid}),
	.s_lval_axis_tready({SUB_54_out_INT_55_2_tready}),
	//rval input
	.s_rval_axis_tdata({select_result_77_tdata}),
	.s_rval_axis_tvalid({select_result_77_tvalid}),
	.s_rval_axis_tready({select_result_77_tready}),
	//output val
	.m_val_axis_tdata({ADD_79_out_INT_80_tdata}),
	.m_val_axis_tvalid({ADD_79_out_INT_80_tvalid}),
	.m_val_axis_tready({ADD_79_out_INT_80_tready})
);

//Arithmetic OP Out
 wire [32-1:0] SUB_81_out_INT_82_tdata;
 wire  SUB_81_out_INT_82_tvalid;
 wire  SUB_81_out_INT_82_tready;

//Arithmetic OP Out
 wire [32-1:0] SUB_81_out_INT_82_0_tdata;
 wire  SUB_81_out_INT_82_0_tvalid;
 wire  SUB_81_out_INT_82_0_tready;

//Arithmetic OP Out
 wire [32-1:0] SUB_81_out_INT_82_1_tdata;
 wire  SUB_81_out_INT_82_1_tvalid;
 wire  SUB_81_out_INT_82_1_tready;

//Arithmetic OP Out
 wire [32-1:0] SUB_81_out_INT_82_2_tdata;
 wire  SUB_81_out_INT_82_2_tvalid;
 wire  SUB_81_out_INT_82_2_tready;

//Arithmetic OP Out
 wire [32-1:0] SUB_81_out_INT_82_3_tdata;
 wire  SUB_81_out_INT_82_3_tvalid;
 wire  SUB_81_out_INT_82_3_tready;

//Arithmetic OP Out
 wire [32-1:0] SUB_81_out_INT_82_4_tdata;
 wire  SUB_81_out_INT_82_4_tvalid;
 wire  SUB_81_out_INT_82_4_tready;

axis_replication#(
.DATA_WIDTH(32),
.IF_STREAM(0),
.REAPLICA_COUNT(5)
)axis_replication_83(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.s_axis_in_tdata({SUB_81_out_INT_82_tdata}),
	.s_axis_in_tvalid({SUB_81_out_INT_82_tvalid}),
	.s_axis_in_tready({SUB_81_out_INT_82_tready}),
	//
	.m_axis_out_tdata({SUB_81_out_INT_82_0_tdata,SUB_81_out_INT_82_1_tdata,SUB_81_out_INT_82_2_tdata,SUB_81_out_INT_82_3_tdata,SUB_81_out_INT_82_4_tdata}),
	.m_axis_out_tvalid({SUB_81_out_INT_82_0_tvalid,SUB_81_out_INT_82_1_tvalid,SUB_81_out_INT_82_2_tvalid,SUB_81_out_INT_82_3_tvalid,SUB_81_out_INT_82_4_tvalid}),
	.m_axis_out_tready({SUB_81_out_INT_82_0_tready,SUB_81_out_INT_82_1_tready,SUB_81_out_INT_82_2_tready,SUB_81_out_INT_82_3_tready,SUB_81_out_INT_82_4_tready})
);

ALU#(
.LVAL_SIZE(32),
.RVAL_SIZE(32),
.RESULT_SIZE(32),
.OPID(0)
)SUB_81(
	 .clk(clk), 
	 .rst(rst) ,
	//lval input
	.s_lval_axis_tdata({struct_accessed_INT_58_2_tdata}),
	.s_lval_axis_tvalid({struct_accessed_INT_58_2_tvalid}),
	.s_lval_axis_tready({struct_accessed_INT_58_2_tready}),
	//rval input
	.s_rval_axis_tdata({ADD_79_out_INT_80_tdata}),
	.s_rval_axis_tvalid({ADD_79_out_INT_80_tvalid}),
	.s_rval_axis_tready({ADD_79_out_INT_80_tready}),
	//output val
	.m_val_axis_tdata({SUB_81_out_INT_82_tdata}),
	.m_val_axis_tvalid({SUB_81_out_INT_82_tvalid}),
	.m_val_axis_tready({SUB_81_out_INT_82_tready})
);

//Arithmetic OP Out
 wire [1-1:0] GT_84_out_INT_85_tdata;
 wire  GT_84_out_INT_85_tvalid;
 wire  GT_84_out_INT_85_tready;

//Arithmetic OP Out
 wire [1-1:0] GT_84_out_INT_85_0_tdata;
 wire  GT_84_out_INT_85_0_tvalid;
 wire  GT_84_out_INT_85_0_tready;

//Arithmetic OP Out
 wire [1-1:0] GT_84_out_INT_85_1_tdata;
 wire  GT_84_out_INT_85_1_tvalid;
 wire  GT_84_out_INT_85_1_tready;

axis_replication#(
.DATA_WIDTH(1),
.IF_STREAM(0),
.REAPLICA_COUNT(2)
)axis_replication_86(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.s_axis_in_tdata({GT_84_out_INT_85_tdata}),
	.s_axis_in_tvalid({GT_84_out_INT_85_tvalid}),
	.s_axis_in_tready({GT_84_out_INT_85_tready}),
	//
	.m_axis_out_tdata({GT_84_out_INT_85_0_tdata,GT_84_out_INT_85_1_tdata}),
	.m_axis_out_tvalid({GT_84_out_INT_85_0_tvalid,GT_84_out_INT_85_1_tvalid}),
	.m_axis_out_tready({GT_84_out_INT_85_0_tready,GT_84_out_INT_85_1_tready})
);

ALU#(
.LVAL_SIZE(32),
.RVAL_SIZE(64),
.RESULT_SIZE(1),
.OPID(4)
)GT_84(
	 .clk(clk), 
	 .rst(rst) ,
	//lval input
	.s_lval_axis_tdata({SUB_81_out_INT_82_0_tdata}),
	.s_lval_axis_tvalid({SUB_81_out_INT_82_0_tvalid}),
	.s_lval_axis_tready({SUB_81_out_INT_82_0_tready}),
	//rval input
	.s_rval_axis_tdata({const_INT_40_tdata}),
	.s_rval_axis_tvalid({const_INT_40_tvalid}),
	.s_rval_axis_tready({const_INT_40_tready}),
	//output val
	.m_val_axis_tdata({GT_84_out_INT_85_tdata}),
	.m_val_axis_tvalid({GT_84_out_INT_85_tvalid}),
	.m_val_axis_tready({GT_84_out_INT_85_tready})
);

//Arithmetic OP Out
 wire [32-1:0] SUB_87_out_INT_88_tdata;
 wire  SUB_87_out_INT_88_tvalid;
 wire  SUB_87_out_INT_88_tready;

ALU#(
.LVAL_SIZE(32),
.RVAL_SIZE(32),
.RESULT_SIZE(32),
.OPID(0)
)SUB_87(
	 .clk(clk), 
	 .rst(rst) ,
	//lval input
	.s_lval_axis_tdata({struct_accessed_INT_64_2_tdata}),
	.s_lval_axis_tvalid({struct_accessed_INT_64_2_tvalid}),
	.s_lval_axis_tready({struct_accessed_INT_64_2_tready}),
	//rval input
	.s_rval_axis_tdata({SUB_81_out_INT_82_1_tdata}),
	.s_rval_axis_tvalid({SUB_81_out_INT_82_1_tvalid}),
	.s_rval_axis_tready({SUB_81_out_INT_82_1_tready}),
	//output val
	.m_val_axis_tdata({SUB_87_out_INT_88_tdata}),
	.m_val_axis_tvalid({SUB_87_out_INT_88_tvalid}),
	.m_val_axis_tready({SUB_87_out_INT_88_tready})
);

//struct_assign_89 output struct
 wire [64-1:0] structvar_90_tdata;
 wire  structvar_90_tvalid;
 wire  structvar_90_tready;

struct_assign#(
.STRUCT_WIDTH(64),
.ASSIGN_OFFSET(32),
.ASSIGN_SIZE(32)
)struct_assign_89(
	 .clk(clk), 
	 .rst(rst) ,
	//input struct
	.s_struct_axis_tdata({structvar_76_tdata}),
	.s_struct_axis_tvalid({structvar_76_tvalid}),
	.s_struct_axis_tready({structvar_76_tready}),
	//input val
	.s_assignv_axis_tdata({SUB_81_out_INT_82_2_tdata}),
	.s_assignv_axis_tvalid({SUB_81_out_INT_82_2_tvalid}),
	.s_assignv_axis_tready({SUB_81_out_INT_82_2_tready}),
	//output struct
	.m_struct_axis_tdata({structvar_90_tdata}),
	.m_struct_axis_tvalid({structvar_90_tvalid}),
	.m_struct_axis_tready({structvar_90_tready})
);

//struct_assign_91 output struct
 wire [256-1:0] structvar_92_tdata;
 wire  structvar_92_tvalid;
 wire  structvar_92_tready;

//struct_assign_91 output struct
 wire [256-1:0] structvar_92_0_tdata;
 wire  structvar_92_0_tvalid;
 wire  structvar_92_0_tready;

//struct_assign_91 output struct
 wire [256-1:0] structvar_92_1_tdata;
 wire  structvar_92_1_tvalid;
 wire  structvar_92_1_tready;

axis_replication#(
.DATA_WIDTH(256),
.IF_STREAM(0),
.REAPLICA_COUNT(2)
)axis_replication_93(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.s_axis_in_tdata({structvar_92_tdata}),
	.s_axis_in_tvalid({structvar_92_tvalid}),
	.s_axis_in_tready({structvar_92_tready}),
	//
	.m_axis_out_tdata({structvar_92_0_tdata,structvar_92_1_tdata}),
	.m_axis_out_tvalid({structvar_92_0_tvalid,structvar_92_1_tvalid}),
	.m_axis_out_tready({structvar_92_0_tready,structvar_92_1_tready})
);

struct_assign#(
.STRUCT_WIDTH(256),
.ASSIGN_OFFSET(96),
.ASSIGN_SIZE(32)
)struct_assign_91(
	 .clk(clk), 
	 .rst(rst) ,
	//input struct
	.s_struct_axis_tdata({lookedup_STRUCT_46_3_tdata}),
	.s_struct_axis_tvalid({lookedup_STRUCT_46_3_tvalid}),
	.s_struct_axis_tready({lookedup_STRUCT_46_3_tready}),
	//input val
	.s_assignv_axis_tdata({SUB_87_out_INT_88_tdata}),
	.s_assignv_axis_tvalid({SUB_87_out_INT_88_tvalid}),
	.s_assignv_axis_tready({SUB_87_out_INT_88_tready}),
	//output struct
	.m_struct_axis_tdata({structvar_92_tdata}),
	.m_struct_axis_tvalid({structvar_92_tvalid}),
	.m_struct_axis_tready({structvar_92_tready})
);

//Access Struct
 wire [32-1:0] struct_accessed_INT_95_tdata;
 wire  struct_accessed_INT_95_tvalid;
 wire  struct_accessed_INT_95_tready;

struct_access#(
.STRUCT_WIDTH(256),
.ACCESS_OFFSET(128),
.ACCESS_SIZE(32)
)struct_access_94(
	 .clk(clk), 
	 .rst(rst) ,
	//struct input
	.s_struct_axis_tdata({structvar_92_0_tdata}),
	.s_struct_axis_tvalid({structvar_92_0_tvalid}),
	.s_struct_axis_tready({structvar_92_0_tready}),
	//output val
	.m_val_axis_tdata({struct_accessed_INT_95_tdata}),
	.m_val_axis_tvalid({struct_accessed_INT_95_tvalid}),
	.m_val_axis_tready({struct_accessed_INT_95_tready})
);

//replicated guard condition
 wire [1-1:0] replicated_guard_cond_96_tdata;
 wire  replicated_guard_cond_96_tvalid;
 wire  replicated_guard_cond_96_tready;

//replicated guard condition
 wire [1-1:0] replicated_guard_cond_97_tdata;
 wire  replicated_guard_cond_97_tvalid;
 wire  replicated_guard_cond_97_tready;

//replicated guard condition
 wire [1-1:0] replicated_guard_cond_98_tdata;
 wire  replicated_guard_cond_98_tvalid;
 wire  replicated_guard_cond_98_tready;

//replicated guard condition
 wire [1-1:0] replicated_guard_cond_99_tdata;
 wire  replicated_guard_cond_99_tvalid;
 wire  replicated_guard_cond_99_tready;

//replicated guard condition
 wire [1-1:0] replicated_guard_cond_100_tdata;
 wire  replicated_guard_cond_100_tvalid;
 wire  replicated_guard_cond_100_tready;

//replicated guard condition
 wire [1-1:0] replicated_guard_cond_101_tdata;
 wire  replicated_guard_cond_101_tvalid;
 wire  replicated_guard_cond_101_tready;

guard_pred#(
.COND_WIDTH(2),
.REPLICATED_OUT_NUM(6),
.GROUND_TRUTH(3)
)guard_pred_102(
	 .clk(clk), 
	 .rst(rst) ,
	//guard condition
	.s_guard_cond_tdata({GT_84_out_INT_85_0_tdata,LE_70_out_INT_71_0_tdata}),
	.s_guard_cond_tvalid({GT_84_out_INT_85_0_tvalid,LE_70_out_INT_71_0_tvalid}),
	.s_guard_cond_tready({GT_84_out_INT_85_0_tready,LE_70_out_INT_71_0_tready}),
	//replicated guard condition
	.m_guard_cond_tdata({replicated_guard_cond_96_tdata,replicated_guard_cond_97_tdata,replicated_guard_cond_98_tdata,replicated_guard_cond_99_tdata,replicated_guard_cond_100_tdata,replicated_guard_cond_101_tdata}),
	.m_guard_cond_tvalid({replicated_guard_cond_96_tvalid,replicated_guard_cond_97_tvalid,replicated_guard_cond_98_tvalid,replicated_guard_cond_99_tvalid,replicated_guard_cond_100_tvalid,replicated_guard_cond_101_tvalid}),
	.m_guard_cond_tready({replicated_guard_cond_96_tready,replicated_guard_cond_97_tready,replicated_guard_cond_98_tready,replicated_guard_cond_99_tready,replicated_guard_cond_100_tready,replicated_guard_cond_101_tready})
);

//Outport Assign Src Value-- guarded
 wire [512-1:0] arg_29_0_guarded_tdata;
 wire [64-1:0] arg_29_0_guarded_tkeep;
 wire  arg_29_0_guarded_tvalid;
 wire  arg_29_0_guarded_tready;
 wire  arg_29_0_guarded_tlast;

guard#(
.DATA_WIDTH(512),
.IF_STREAM(1)
)guard_103(
	 .clk(clk), 
	 .rst(rst) ,
	//input val
	.s_guard_axis_tdata({arg_29_0_tdata}),
	.s_guard_axis_tkeep({arg_29_0_tkeep}),
	.s_guard_axis_tlast({arg_29_0_tlast}),
	.s_guard_axis_tvalid({arg_29_0_tvalid}),
	.s_guard_axis_tready({arg_29_0_tready}),
	//output val
	.m_guard_axis_tdata({arg_29_0_guarded_tdata}),
	.m_guard_axis_tkeep({arg_29_0_guarded_tkeep}),
	.m_guard_axis_tlast({arg_29_0_guarded_tlast}),
	.m_guard_axis_tvalid({arg_29_0_guarded_tvalid}),
	.m_guard_axis_tready({arg_29_0_guarded_tready}),
	//guard condition
	.s_guard_cond_tdata({replicated_guard_cond_96_tdata}),
	.s_guard_cond_tvalid({replicated_guard_cond_96_tvalid}),
	.s_guard_cond_tready({replicated_guard_cond_96_tready})
);

 assign DMA_WRITE_1_tdata = arg_29_0_guarded_tdata;
 assign DMA_WRITE_1_tvalid = arg_29_0_guarded_tvalid;
 assign arg_29_0_guarded_tready = DMA_WRITE_1_tready;
 assign DMA_WRITE_1_tkeep = arg_29_0_guarded_tkeep;
 assign DMA_WRITE_1_tlast = arg_29_0_guarded_tlast;

//Outport Assign Src Value-- guarded
 wire [64-1:0] structvar_90_guarded_tdata;
 wire  structvar_90_guarded_tvalid;
 wire  structvar_90_guarded_tready;

guard#(
.DATA_WIDTH(64),
.IF_STREAM(0)
)guard_104(
	 .clk(clk), 
	 .rst(rst) ,
	//input val
	.s_guard_axis_tdata({structvar_90_tdata}),
	.s_guard_axis_tvalid({structvar_90_tvalid}),
	.s_guard_axis_tready({structvar_90_tready}),
	//output val
	.m_guard_axis_tdata({structvar_90_guarded_tdata}),
	.m_guard_axis_tvalid({structvar_90_guarded_tvalid}),
	.m_guard_axis_tready({structvar_90_guarded_tready}),
	//guard condition
	.s_guard_cond_tdata({replicated_guard_cond_97_tdata}),
	.s_guard_cond_tvalid({replicated_guard_cond_97_tvalid}),
	.s_guard_cond_tready({replicated_guard_cond_97_tready})
);

 assign DMA_WRITE_2_tdata = structvar_90_guarded_tdata;
 assign DMA_WRITE_2_tvalid = structvar_90_guarded_tvalid;
 assign structvar_90_guarded_tready = DMA_WRITE_2_tready;

//Outport Assign Src Value-- guarded
 wire [512-1:0] arg_29_1_guarded_tdata;
 wire [64-1:0] arg_29_1_guarded_tkeep;
 wire  arg_29_1_guarded_tvalid;
 wire  arg_29_1_guarded_tready;
 wire  arg_29_1_guarded_tlast;

guard#(
.DATA_WIDTH(512),
.IF_STREAM(1)
)guard_105(
	 .clk(clk), 
	 .rst(rst) ,
	//input val
	.s_guard_axis_tdata({arg_29_1_tdata}),
	.s_guard_axis_tkeep({arg_29_1_tkeep}),
	.s_guard_axis_tlast({arg_29_1_tlast}),
	.s_guard_axis_tvalid({arg_29_1_tvalid}),
	.s_guard_axis_tready({arg_29_1_tready}),
	//output val
	.m_guard_axis_tdata({arg_29_1_guarded_tdata}),
	.m_guard_axis_tkeep({arg_29_1_guarded_tkeep}),
	.m_guard_axis_tlast({arg_29_1_guarded_tlast}),
	.m_guard_axis_tvalid({arg_29_1_guarded_tvalid}),
	.m_guard_axis_tready({arg_29_1_guarded_tready}),
	//guard condition
	.s_guard_cond_tdata({replicated_guard_cond_98_tdata}),
	.s_guard_cond_tvalid({replicated_guard_cond_98_tvalid}),
	.s_guard_cond_tready({replicated_guard_cond_98_tready})
);

 assign DMA_WRITE_3_tdata = arg_29_1_guarded_tdata;
 assign DMA_WRITE_3_tvalid = arg_29_1_guarded_tvalid;
 assign arg_29_1_guarded_tready = DMA_WRITE_3_tready;
 assign DMA_WRITE_3_tkeep = arg_29_1_guarded_tkeep;
 assign DMA_WRITE_3_tlast = arg_29_1_guarded_tlast;

//Outport Assign Src Value-- guarded
 wire [184-1:0] arg_30_0_guarded_tdata;
 wire  arg_30_0_guarded_tvalid;
 wire  arg_30_0_guarded_tready;

guard#(
.DATA_WIDTH(184),
.IF_STREAM(0)
)guard_106(
	 .clk(clk), 
	 .rst(rst) ,
	//input val
	.s_guard_axis_tdata({arg_30_0_tdata}),
	.s_guard_axis_tvalid({arg_30_0_tvalid}),
	.s_guard_axis_tready({arg_30_0_tready}),
	//output val
	.m_guard_axis_tdata({arg_30_0_guarded_tdata}),
	.m_guard_axis_tvalid({arg_30_0_guarded_tvalid}),
	.m_guard_axis_tready({arg_30_0_guarded_tready}),
	//guard condition
	.s_guard_cond_tdata({replicated_guard_cond_99_tdata}),
	.s_guard_cond_tvalid({replicated_guard_cond_99_tvalid}),
	.s_guard_cond_tready({replicated_guard_cond_99_tready})
);

 assign DMA_WRITE_4_tdata = arg_30_0_guarded_tdata;
 assign DMA_WRITE_4_tvalid = arg_30_0_guarded_tvalid;
 assign arg_30_0_guarded_tready = DMA_WRITE_4_tready;

//Outport Assign Src Value-- guarded
 wire [112-1:0] arg_31_0_guarded_tdata;
 wire  arg_31_0_guarded_tvalid;
 wire  arg_31_0_guarded_tready;

guard#(
.DATA_WIDTH(112),
.IF_STREAM(0)
)guard_107(
	 .clk(clk), 
	 .rst(rst) ,
	//input val
	.s_guard_axis_tdata({arg_31_0_tdata}),
	.s_guard_axis_tvalid({arg_31_0_tvalid}),
	.s_guard_axis_tready({arg_31_0_tready}),
	//output val
	.m_guard_axis_tdata({arg_31_0_guarded_tdata}),
	.m_guard_axis_tvalid({arg_31_0_guarded_tvalid}),
	.m_guard_axis_tready({arg_31_0_guarded_tready}),
	//guard condition
	.s_guard_cond_tdata({replicated_guard_cond_100_tdata}),
	.s_guard_cond_tvalid({replicated_guard_cond_100_tvalid}),
	.s_guard_cond_tready({replicated_guard_cond_100_tready})
);

 assign DMA_WRITE_5_tdata = arg_31_0_guarded_tdata;
 assign DMA_WRITE_5_tvalid = arg_31_0_guarded_tvalid;
 assign arg_31_0_guarded_tready = DMA_WRITE_5_tready;

//Outport Assign Src Value-- guarded
 wire [160-1:0] arg_32_0_guarded_tdata;
 wire  arg_32_0_guarded_tvalid;
 wire  arg_32_0_guarded_tready;

guard#(
.DATA_WIDTH(160),
.IF_STREAM(0)
)guard_108(
	 .clk(clk), 
	 .rst(rst) ,
	//input val
	.s_guard_axis_tdata({arg_32_0_tdata}),
	.s_guard_axis_tvalid({arg_32_0_tvalid}),
	.s_guard_axis_tready({arg_32_0_tready}),
	//output val
	.m_guard_axis_tdata({arg_32_0_guarded_tdata}),
	.m_guard_axis_tvalid({arg_32_0_guarded_tvalid}),
	.m_guard_axis_tready({arg_32_0_guarded_tready}),
	//guard condition
	.s_guard_cond_tdata({replicated_guard_cond_101_tdata}),
	.s_guard_cond_tvalid({replicated_guard_cond_101_tvalid}),
	.s_guard_cond_tready({replicated_guard_cond_101_tready})
);

 assign DMA_WRITE_6_tdata = arg_32_0_guarded_tdata;
 assign DMA_WRITE_6_tvalid = arg_32_0_guarded_tvalid;
 assign arg_32_0_guarded_tready = DMA_WRITE_6_tready;

//Arithmetic OP Out
 wire [32-1:0] ADD_109_out_INT_110_tdata;
 wire  ADD_109_out_INT_110_tvalid;
 wire  ADD_109_out_INT_110_tready;

ALU#(
.LVAL_SIZE(32),
.RVAL_SIZE(32),
.RESULT_SIZE(32),
.OPID(1)
)ADD_109(
	 .clk(clk), 
	 .rst(rst) ,
	//lval input
	.s_lval_axis_tdata({struct_accessed_INT_95_tdata}),
	.s_lval_axis_tvalid({struct_accessed_INT_95_tvalid}),
	.s_lval_axis_tready({struct_accessed_INT_95_tready}),
	//rval input
	.s_rval_axis_tdata({SUB_81_out_INT_82_3_tdata}),
	.s_rval_axis_tvalid({SUB_81_out_INT_82_3_tvalid}),
	.s_rval_axis_tready({SUB_81_out_INT_82_3_tready}),
	//output val
	.m_val_axis_tdata({ADD_109_out_INT_110_tdata}),
	.m_val_axis_tvalid({ADD_109_out_INT_110_tvalid}),
	.m_val_axis_tready({ADD_109_out_INT_110_tready})
);

//struct_assign_111 output struct
 wire [256-1:0] structvar_112_tdata;
 wire  structvar_112_tvalid;
 wire  structvar_112_tready;

//struct_assign_111 output struct
 wire [256-1:0] structvar_112_0_tdata;
 wire  structvar_112_0_tvalid;
 wire  structvar_112_0_tready;

//struct_assign_111 output struct
 wire [256-1:0] structvar_112_1_tdata;
 wire  structvar_112_1_tvalid;
 wire  structvar_112_1_tready;

axis_replication#(
.DATA_WIDTH(256),
.IF_STREAM(0),
.REAPLICA_COUNT(2)
)axis_replication_113(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.s_axis_in_tdata({structvar_112_tdata}),
	.s_axis_in_tvalid({structvar_112_tvalid}),
	.s_axis_in_tready({structvar_112_tready}),
	//
	.m_axis_out_tdata({structvar_112_0_tdata,structvar_112_1_tdata}),
	.m_axis_out_tvalid({structvar_112_0_tvalid,structvar_112_1_tvalid}),
	.m_axis_out_tready({structvar_112_0_tready,structvar_112_1_tready})
);

struct_assign#(
.STRUCT_WIDTH(256),
.ASSIGN_OFFSET(128),
.ASSIGN_SIZE(32)
)struct_assign_111(
	 .clk(clk), 
	 .rst(rst) ,
	//input struct
	.s_struct_axis_tdata({structvar_92_1_tdata}),
	.s_struct_axis_tvalid({structvar_92_1_tvalid}),
	.s_struct_axis_tready({structvar_92_1_tready}),
	//input val
	.s_assignv_axis_tdata({ADD_109_out_INT_110_tdata}),
	.s_assignv_axis_tvalid({ADD_109_out_INT_110_tvalid}),
	.s_assignv_axis_tready({ADD_109_out_INT_110_tready}),
	//output struct
	.m_struct_axis_tdata({structvar_112_tdata}),
	.m_struct_axis_tvalid({structvar_112_tvalid}),
	.m_struct_axis_tready({structvar_112_tready})
);

//Access Struct
 wire [32-1:0] struct_accessed_INT_115_tdata;
 wire  struct_accessed_INT_115_tvalid;
 wire  struct_accessed_INT_115_tready;

struct_access#(
.STRUCT_WIDTH(256),
.ACCESS_OFFSET(160),
.ACCESS_SIZE(32)
)struct_access_114(
	 .clk(clk), 
	 .rst(rst) ,
	//struct input
	.s_struct_axis_tdata({structvar_112_0_tdata}),
	.s_struct_axis_tvalid({structvar_112_0_tvalid}),
	.s_struct_axis_tready({structvar_112_0_tready}),
	//output val
	.m_val_axis_tdata({struct_accessed_INT_115_tdata}),
	.m_val_axis_tvalid({struct_accessed_INT_115_tvalid}),
	.m_val_axis_tready({struct_accessed_INT_115_tready})
);

//Arithmetic OP Out
 wire [32-1:0] ADD_116_out_INT_117_tdata;
 wire  ADD_116_out_INT_117_tvalid;
 wire  ADD_116_out_INT_117_tready;

ALU#(
.LVAL_SIZE(32),
.RVAL_SIZE(32),
.RESULT_SIZE(32),
.OPID(1)
)ADD_116(
	 .clk(clk), 
	 .rst(rst) ,
	//lval input
	.s_lval_axis_tdata({struct_accessed_INT_115_tdata}),
	.s_lval_axis_tvalid({struct_accessed_INT_115_tvalid}),
	.s_lval_axis_tready({struct_accessed_INT_115_tready}),
	//rval input
	.s_rval_axis_tdata({SUB_81_out_INT_82_4_tdata}),
	.s_rval_axis_tvalid({SUB_81_out_INT_82_4_tvalid}),
	.s_rval_axis_tready({SUB_81_out_INT_82_4_tready}),
	//output val
	.m_val_axis_tdata({ADD_116_out_INT_117_tdata}),
	.m_val_axis_tvalid({ADD_116_out_INT_117_tvalid}),
	.m_val_axis_tready({ADD_116_out_INT_117_tready})
);

//struct_assign_118 output struct
 wire [256-1:0] structvar_119_tdata;
 wire  structvar_119_tvalid;
 wire  structvar_119_tready;

struct_assign#(
.STRUCT_WIDTH(256),
.ASSIGN_OFFSET(160),
.ASSIGN_SIZE(32)
)struct_assign_118(
	 .clk(clk), 
	 .rst(rst) ,
	//input struct
	.s_struct_axis_tdata({structvar_112_1_tdata}),
	.s_struct_axis_tvalid({structvar_112_1_tvalid}),
	.s_struct_axis_tready({structvar_112_1_tready}),
	//input val
	.s_assignv_axis_tdata({ADD_116_out_INT_117_tdata}),
	.s_assignv_axis_tvalid({ADD_116_out_INT_117_tvalid}),
	.s_assignv_axis_tready({ADD_116_out_INT_117_tready}),
	//output struct
	.m_struct_axis_tdata({structvar_119_tdata}),
	.m_struct_axis_tvalid({structvar_119_tvalid}),
	.m_struct_axis_tready({structvar_119_tready})
);

//
 wire [256-1:0] select_result_120_tdata;
 wire  select_result_120_tvalid;
 wire  select_result_120_tready;

//
 wire [256-1:0] select_result_120_0_tdata;
 wire  select_result_120_0_tvalid;
 wire  select_result_120_0_tready;

//
 wire [256-1:0] select_result_120_1_tdata;
 wire  select_result_120_1_tvalid;
 wire  select_result_120_1_tready;

//
 wire [256-1:0] select_result_120_2_tdata;
 wire  select_result_120_2_tvalid;
 wire  select_result_120_2_tready;

//
 wire [256-1:0] select_result_120_3_tdata;
 wire  select_result_120_3_tvalid;
 wire  select_result_120_3_tready;

axis_replication#(
.DATA_WIDTH(256),
.IF_STREAM(0),
.REAPLICA_COUNT(4)
)axis_replication_121(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.s_axis_in_tdata({select_result_120_tdata}),
	.s_axis_in_tvalid({select_result_120_tvalid}),
	.s_axis_in_tready({select_result_120_tready}),
	//
	.m_axis_out_tdata({select_result_120_0_tdata,select_result_120_1_tdata,select_result_120_2_tdata,select_result_120_3_tdata}),
	.m_axis_out_tvalid({select_result_120_0_tvalid,select_result_120_1_tvalid,select_result_120_2_tvalid,select_result_120_3_tvalid}),
	.m_axis_out_tready({select_result_120_0_tready,select_result_120_1_tready,select_result_120_2_tready,select_result_120_3_tready})
);

select#(
.VAL_WIDTH(256),
.COND_WIDTH(1)
)select_122(
	 .clk(clk), 
	 .rst(rst) ,
	//select condition
	.s_cond_axis_tdata({GT_84_out_INT_85_1_tdata}),
	.s_cond_axis_tvalid({GT_84_out_INT_85_1_tvalid}),
	.s_cond_axis_tready({GT_84_out_INT_85_1_tready}),
	//select true val
	.s_true_val_axis_tdata({structvar_119_tdata}),
	.s_true_val_axis_tvalid({structvar_119_tvalid}),
	.s_true_val_axis_tready({structvar_119_tready}),
	//select false val
	.s_false_val_axis_tdata({lookedup_STRUCT_46_4_tdata}),
	.s_false_val_axis_tvalid({lookedup_STRUCT_46_4_tvalid}),
	.s_false_val_axis_tready({lookedup_STRUCT_46_4_tready}),
	//select result
	.m_val_axis_tdata({select_result_120_tdata}),
	.m_val_axis_tvalid({select_result_120_tvalid}),
	.m_val_axis_tready({select_result_120_tready})
);

//replicated guard condition
 wire [1-1:0] replicated_guard_cond_123_tdata;
 wire  replicated_guard_cond_123_tvalid;
 wire  replicated_guard_cond_123_tready;

//replicated guard condition
 wire [1-1:0] replicated_guard_cond_124_tdata;
 wire  replicated_guard_cond_124_tvalid;
 wire  replicated_guard_cond_124_tready;

guard_pred#(
.COND_WIDTH(1),
.REPLICATED_OUT_NUM(2),
.GROUND_TRUTH(1)
)guard_pred_125(
	 .clk(clk), 
	 .rst(rst) ,
	//guard condition
	.s_guard_cond_tdata({LE_70_out_INT_71_1_tdata}),
	.s_guard_cond_tvalid({LE_70_out_INT_71_1_tvalid}),
	.s_guard_cond_tready({LE_70_out_INT_71_1_tready}),
	//replicated guard condition
	.m_guard_cond_tdata({replicated_guard_cond_123_tdata,replicated_guard_cond_124_tdata}),
	.m_guard_cond_tvalid({replicated_guard_cond_123_tvalid,replicated_guard_cond_124_tvalid}),
	.m_guard_cond_tready({replicated_guard_cond_123_tready,replicated_guard_cond_124_tready})
);

//-- guarded
 wire [16-1:0] bitcasted_44_1_guarded_tdata;
 wire  bitcasted_44_1_guarded_tvalid;
 wire  bitcasted_44_1_guarded_tready;

guard#(
.DATA_WIDTH(16),
.IF_STREAM(0)
)guard_126(
	 .clk(clk), 
	 .rst(rst) ,
	//input val
	.s_guard_axis_tdata({bitcasted_44_1_tdata}),
	.s_guard_axis_tvalid({bitcasted_44_1_tvalid}),
	.s_guard_axis_tready({bitcasted_44_1_tready}),
	//output val
	.m_guard_axis_tdata({bitcasted_44_1_guarded_tdata}),
	.m_guard_axis_tvalid({bitcasted_44_1_guarded_tvalid}),
	.m_guard_axis_tready({bitcasted_44_1_guarded_tready}),
	//guard condition
	.s_guard_cond_tdata({replicated_guard_cond_123_tdata}),
	.s_guard_cond_tvalid({replicated_guard_cond_123_tvalid}),
	.s_guard_cond_tready({replicated_guard_cond_123_tready})
);

//-- guarded
 wire [256-1:0] select_result_120_0_guarded_tdata;
 wire  select_result_120_0_guarded_tvalid;
 wire  select_result_120_0_guarded_tready;

guard#(
.DATA_WIDTH(256),
.IF_STREAM(0)
)guard_127(
	 .clk(clk), 
	 .rst(rst) ,
	//input val
	.s_guard_axis_tdata({select_result_120_0_tdata}),
	.s_guard_axis_tvalid({select_result_120_0_tvalid}),
	.s_guard_axis_tready({select_result_120_0_tready}),
	//output val
	.m_guard_axis_tdata({select_result_120_0_guarded_tdata}),
	.m_guard_axis_tvalid({select_result_120_0_guarded_tvalid}),
	.m_guard_axis_tready({select_result_120_0_guarded_tready}),
	//guard condition
	.s_guard_cond_tdata({replicated_guard_cond_124_tdata}),
	.s_guard_cond_tvalid({replicated_guard_cond_124_tvalid}),
	.s_guard_cond_tready({replicated_guard_cond_124_tready})
);

 assign update_p_0_req_index = bitcasted_44_1_guarded_tdata;
 assign update_p_0_req_index_valid = bitcasted_44_1_guarded_tvalid;
 assign bitcasted_44_1_guarded_tready = update_p_0_req_index_ready;

 assign update_p_0_req_data = select_result_120_0_guarded_tdata;
 assign update_p_0_req_data_valid = select_result_120_0_guarded_tvalid;
 assign select_result_120_0_guarded_tready = update_p_0_req_data_ready;

//Access Struct
 wire [32-1:0] struct_accessed_INT_129_tdata;
 wire  struct_accessed_INT_129_tvalid;
 wire  struct_accessed_INT_129_tready;

struct_access#(
.STRUCT_WIDTH(256),
.ACCESS_OFFSET(0),
.ACCESS_SIZE(32)
)struct_access_128(
	 .clk(clk), 
	 .rst(rst) ,
	//struct input
	.s_struct_axis_tdata({select_result_120_1_tdata}),
	.s_struct_axis_tvalid({select_result_120_1_tvalid}),
	.s_struct_axis_tready({select_result_120_1_tready}),
	//output val
	.m_val_axis_tdata({struct_accessed_INT_129_tdata}),
	.m_val_axis_tvalid({struct_accessed_INT_129_tvalid}),
	.m_val_axis_tready({struct_accessed_INT_129_tready})
);

//Access Struct
 wire [32-1:0] struct_accessed_INT_131_tdata;
 wire  struct_accessed_INT_131_tvalid;
 wire  struct_accessed_INT_131_tready;

struct_access#(
.STRUCT_WIDTH(256),
.ACCESS_OFFSET(128),
.ACCESS_SIZE(32)
)struct_access_130(
	 .clk(clk), 
	 .rst(rst) ,
	//struct input
	.s_struct_axis_tdata({select_result_120_2_tdata}),
	.s_struct_axis_tvalid({select_result_120_2_tvalid}),
	.s_struct_axis_tready({select_result_120_2_tready}),
	//output val
	.m_val_axis_tdata({struct_accessed_INT_131_tdata}),
	.m_val_axis_tvalid({struct_accessed_INT_131_tvalid}),
	.m_val_axis_tready({struct_accessed_INT_131_tready})
);

//Access Struct
 wire [32-1:0] struct_accessed_INT_133_tdata;
 wire  struct_accessed_INT_133_tvalid;
 wire  struct_accessed_INT_133_tready;

struct_access#(
.STRUCT_WIDTH(256),
.ACCESS_OFFSET(96),
.ACCESS_SIZE(32)
)struct_access_132(
	 .clk(clk), 
	 .rst(rst) ,
	//struct input
	.s_struct_axis_tdata({select_result_120_3_tdata}),
	.s_struct_axis_tvalid({select_result_120_3_tvalid}),
	.s_struct_axis_tready({select_result_120_3_tready}),
	//output val
	.m_val_axis_tdata({struct_accessed_INT_133_tdata}),
	.m_val_axis_tvalid({struct_accessed_INT_133_tvalid}),
	.m_val_axis_tready({struct_accessed_INT_133_tready})
);

//struct_assign_134 output struct
 wire [96-1:0] structvar_135_tdata;
 wire  structvar_135_tvalid;
 wire  structvar_135_tready;

struct_assign#(
.STRUCT_WIDTH(96),
.ASSIGN_OFFSET(0),
.ASSIGN_SIZE(32)
)struct_assign_134(
	 .clk(clk), 
	 .rst(rst) ,
	//input struct
	.s_struct_axis_tdata({inited_STRUCT_49_tdata}),
	.s_struct_axis_tvalid({inited_STRUCT_49_tvalid}),
	.s_struct_axis_tready({inited_STRUCT_49_tready}),
	//input val
	.s_assignv_axis_tdata({struct_accessed_INT_129_tdata}),
	.s_assignv_axis_tvalid({struct_accessed_INT_129_tvalid}),
	.s_assignv_axis_tready({struct_accessed_INT_129_tready}),
	//output struct
	.m_struct_axis_tdata({structvar_135_tdata}),
	.m_struct_axis_tvalid({structvar_135_tvalid}),
	.m_struct_axis_tready({structvar_135_tready})
);

//struct_assign_136 output struct
 wire [96-1:0] structvar_137_tdata;
 wire  structvar_137_tvalid;
 wire  structvar_137_tready;

struct_assign#(
.STRUCT_WIDTH(96),
.ASSIGN_OFFSET(32),
.ASSIGN_SIZE(32)
)struct_assign_136(
	 .clk(clk), 
	 .rst(rst) ,
	//input struct
	.s_struct_axis_tdata({structvar_135_tdata}),
	.s_struct_axis_tvalid({structvar_135_tvalid}),
	.s_struct_axis_tready({structvar_135_tready}),
	//input val
	.s_assignv_axis_tdata({struct_accessed_INT_131_tdata}),
	.s_assignv_axis_tvalid({struct_accessed_INT_131_tvalid}),
	.s_assignv_axis_tready({struct_accessed_INT_131_tready}),
	//output struct
	.m_struct_axis_tdata({structvar_137_tdata}),
	.m_struct_axis_tvalid({structvar_137_tvalid}),
	.m_struct_axis_tready({structvar_137_tready})
);

//struct_assign_138 output struct
 wire [96-1:0] structvar_139_tdata;
 wire  structvar_139_tvalid;
 wire  structvar_139_tready;

struct_assign#(
.STRUCT_WIDTH(96),
.ASSIGN_OFFSET(64),
.ASSIGN_SIZE(32)
)struct_assign_138(
	 .clk(clk), 
	 .rst(rst) ,
	//input struct
	.s_struct_axis_tdata({structvar_137_tdata}),
	.s_struct_axis_tvalid({structvar_137_tvalid}),
	.s_struct_axis_tready({structvar_137_tready}),
	//input val
	.s_assignv_axis_tdata({struct_accessed_INT_133_tdata}),
	.s_assignv_axis_tvalid({struct_accessed_INT_133_tvalid}),
	.s_assignv_axis_tready({struct_accessed_INT_133_tready}),
	//output struct
	.m_struct_axis_tdata({structvar_139_tdata}),
	.m_struct_axis_tvalid({structvar_139_tvalid}),
	.m_struct_axis_tready({structvar_139_tready})
);

//replicated guard condition
 wire [1-1:0] replicated_guard_cond_140_tdata;
 wire  replicated_guard_cond_140_tvalid;
 wire  replicated_guard_cond_140_tready;

//replicated guard condition
 wire [1-1:0] replicated_guard_cond_141_tdata;
 wire  replicated_guard_cond_141_tvalid;
 wire  replicated_guard_cond_141_tready;

//replicated guard condition
 wire [1-1:0] replicated_guard_cond_142_tdata;
 wire  replicated_guard_cond_142_tvalid;
 wire  replicated_guard_cond_142_tready;

//replicated guard condition
 wire [1-1:0] replicated_guard_cond_143_tdata;
 wire  replicated_guard_cond_143_tvalid;
 wire  replicated_guard_cond_143_tready;

//replicated guard condition
 wire [1-1:0] replicated_guard_cond_144_tdata;
 wire  replicated_guard_cond_144_tvalid;
 wire  replicated_guard_cond_144_tready;

guard_pred#(
.COND_WIDTH(1),
.REPLICATED_OUT_NUM(5),
.GROUND_TRUTH(1)
)guard_pred_145(
	 .clk(clk), 
	 .rst(rst) ,
	//guard condition
	.s_guard_cond_tdata({LE_70_out_INT_71_2_tdata}),
	.s_guard_cond_tvalid({LE_70_out_INT_71_2_tvalid}),
	.s_guard_cond_tready({LE_70_out_INT_71_2_tready}),
	//replicated guard condition
	.m_guard_cond_tdata({replicated_guard_cond_140_tdata,replicated_guard_cond_141_tdata,replicated_guard_cond_142_tdata,replicated_guard_cond_143_tdata,replicated_guard_cond_144_tdata}),
	.m_guard_cond_tvalid({replicated_guard_cond_140_tvalid,replicated_guard_cond_141_tvalid,replicated_guard_cond_142_tvalid,replicated_guard_cond_143_tvalid,replicated_guard_cond_144_tvalid}),
	.m_guard_cond_tready({replicated_guard_cond_140_tready,replicated_guard_cond_141_tready,replicated_guard_cond_142_tready,replicated_guard_cond_143_tready,replicated_guard_cond_144_tready})
);

//Outport Assign Src Value-- guarded
 wire [96-1:0] structvar_139_guarded_tdata;
 wire  structvar_139_guarded_tvalid;
 wire  structvar_139_guarded_tready;

guard#(
.DATA_WIDTH(96),
.IF_STREAM(0)
)guard_146(
	 .clk(clk), 
	 .rst(rst) ,
	//input val
	.s_guard_axis_tdata({structvar_139_tdata}),
	.s_guard_axis_tvalid({structvar_139_tvalid}),
	.s_guard_axis_tready({structvar_139_tready}),
	//output val
	.m_guard_axis_tdata({structvar_139_guarded_tdata}),
	.m_guard_axis_tvalid({structvar_139_guarded_tvalid}),
	.m_guard_axis_tready({structvar_139_guarded_tready}),
	//guard condition
	.s_guard_cond_tdata({replicated_guard_cond_140_tdata}),
	.s_guard_cond_tvalid({replicated_guard_cond_140_tvalid}),
	.s_guard_cond_tready({replicated_guard_cond_140_tready})
);

 assign outport_33_1_tdata = structvar_139_guarded_tdata;
 assign outport_33_1_tvalid = structvar_139_guarded_tvalid;
 assign structvar_139_guarded_tready = outport_33_1_tready;

//Outport Assign Src Value-- guarded
 wire [512-1:0] arg_29_2_guarded_tdata;
 wire [64-1:0] arg_29_2_guarded_tkeep;
 wire  arg_29_2_guarded_tvalid;
 wire  arg_29_2_guarded_tready;
 wire  arg_29_2_guarded_tlast;

guard#(
.DATA_WIDTH(512),
.IF_STREAM(1)
)guard_147(
	 .clk(clk), 
	 .rst(rst) ,
	//input val
	.s_guard_axis_tdata({arg_29_2_tdata}),
	.s_guard_axis_tkeep({arg_29_2_tkeep}),
	.s_guard_axis_tlast({arg_29_2_tlast}),
	.s_guard_axis_tvalid({arg_29_2_tvalid}),
	.s_guard_axis_tready({arg_29_2_tready}),
	//output val
	.m_guard_axis_tdata({arg_29_2_guarded_tdata}),
	.m_guard_axis_tkeep({arg_29_2_guarded_tkeep}),
	.m_guard_axis_tlast({arg_29_2_guarded_tlast}),
	.m_guard_axis_tvalid({arg_29_2_guarded_tvalid}),
	.m_guard_axis_tready({arg_29_2_guarded_tready}),
	//guard condition
	.s_guard_cond_tdata({replicated_guard_cond_141_tdata}),
	.s_guard_cond_tvalid({replicated_guard_cond_141_tvalid}),
	.s_guard_cond_tready({replicated_guard_cond_141_tready})
);

 assign outport_33_2_tdata = arg_29_2_guarded_tdata;
 assign outport_33_2_tvalid = arg_29_2_guarded_tvalid;
 assign arg_29_2_guarded_tready = outport_33_2_tready;
 assign outport_33_2_tkeep = arg_29_2_guarded_tkeep;
 assign outport_33_2_tlast = arg_29_2_guarded_tlast;

//Outport Assign Src Value-- guarded
 wire [184-1:0] arg_30_1_guarded_tdata;
 wire  arg_30_1_guarded_tvalid;
 wire  arg_30_1_guarded_tready;

guard#(
.DATA_WIDTH(184),
.IF_STREAM(0)
)guard_148(
	 .clk(clk), 
	 .rst(rst) ,
	//input val
	.s_guard_axis_tdata({arg_30_1_tdata}),
	.s_guard_axis_tvalid({arg_30_1_tvalid}),
	.s_guard_axis_tready({arg_30_1_tready}),
	//output val
	.m_guard_axis_tdata({arg_30_1_guarded_tdata}),
	.m_guard_axis_tvalid({arg_30_1_guarded_tvalid}),
	.m_guard_axis_tready({arg_30_1_guarded_tready}),
	//guard condition
	.s_guard_cond_tdata({replicated_guard_cond_142_tdata}),
	.s_guard_cond_tvalid({replicated_guard_cond_142_tvalid}),
	.s_guard_cond_tready({replicated_guard_cond_142_tready})
);

 assign outport_33_3_tdata = arg_30_1_guarded_tdata;
 assign outport_33_3_tvalid = arg_30_1_guarded_tvalid;
 assign arg_30_1_guarded_tready = outport_33_3_tready;

//Outport Assign Src Value-- guarded
 wire [112-1:0] arg_31_1_guarded_tdata;
 wire  arg_31_1_guarded_tvalid;
 wire  arg_31_1_guarded_tready;

guard#(
.DATA_WIDTH(112),
.IF_STREAM(0)
)guard_149(
	 .clk(clk), 
	 .rst(rst) ,
	//input val
	.s_guard_axis_tdata({arg_31_1_tdata}),
	.s_guard_axis_tvalid({arg_31_1_tvalid}),
	.s_guard_axis_tready({arg_31_1_tready}),
	//output val
	.m_guard_axis_tdata({arg_31_1_guarded_tdata}),
	.m_guard_axis_tvalid({arg_31_1_guarded_tvalid}),
	.m_guard_axis_tready({arg_31_1_guarded_tready}),
	//guard condition
	.s_guard_cond_tdata({replicated_guard_cond_143_tdata}),
	.s_guard_cond_tvalid({replicated_guard_cond_143_tvalid}),
	.s_guard_cond_tready({replicated_guard_cond_143_tready})
);

 assign outport_33_4_tdata = arg_31_1_guarded_tdata;
 assign outport_33_4_tvalid = arg_31_1_guarded_tvalid;
 assign arg_31_1_guarded_tready = outport_33_4_tready;

//Outport Assign Src Value-- guarded
 wire [160-1:0] arg_32_1_guarded_tdata;
 wire  arg_32_1_guarded_tvalid;
 wire  arg_32_1_guarded_tready;

guard#(
.DATA_WIDTH(160),
.IF_STREAM(0)
)guard_150(
	 .clk(clk), 
	 .rst(rst) ,
	//input val
	.s_guard_axis_tdata({arg_32_1_tdata}),
	.s_guard_axis_tvalid({arg_32_1_tvalid}),
	.s_guard_axis_tready({arg_32_1_tready}),
	//output val
	.m_guard_axis_tdata({arg_32_1_guarded_tdata}),
	.m_guard_axis_tvalid({arg_32_1_guarded_tvalid}),
	.m_guard_axis_tready({arg_32_1_guarded_tready}),
	//guard condition
	.s_guard_cond_tdata({replicated_guard_cond_144_tdata}),
	.s_guard_cond_tvalid({replicated_guard_cond_144_tvalid}),
	.s_guard_cond_tready({replicated_guard_cond_144_tready})
);

 assign outport_33_5_tdata = arg_32_1_guarded_tdata;
 assign outport_33_5_tvalid = arg_32_1_guarded_tvalid;
 assign arg_32_1_guarded_tready = outport_33_5_tready;


endmodule
