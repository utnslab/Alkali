module __handler_OoO_DETECT_OoO_detection#()
(
	 input  wire clk, 
	 input  wire rst,
	//input ports STRUCT
	input wire [96-1:0] arg_28_tdata ,
	input wire  arg_28_tvalid ,
	output wire  arg_28_tready,
	//input ports BUF
	input wire [512-1:0] arg_29_tdata ,
	input wire [64-1:0] arg_29_tkeep ,
	input wire  arg_29_tlast ,
	input wire  arg_29_tvalid ,
	output wire  arg_29_tready,
	//input ports STRUCT
	input wire [184-1:0] arg_30_tdata ,
	input wire  arg_30_tvalid ,
	output wire  arg_30_tready,
	//input ports STRUCT
	input wire [112-1:0] arg_31_tdata ,
	input wire  arg_31_tvalid ,
	output wire  arg_31_tready,
	//input ports STRUCT
	input wire [160-1:0] arg_32_tdata ,
	input wire  arg_32_tvalid ,
	output wire  arg_32_tready,
	//output ports STRUCT
	output wire [96-1:0] outport_33_1_tdata ,
	output wire  outport_33_1_tvalid ,
	input wire  outport_33_1_tready,
	//output ports BUF
	output wire [512-1:0] outport_33_2_tdata ,
	output wire [64-1:0] outport_33_2_tkeep ,
	output wire  outport_33_2_tlast ,
	output wire  outport_33_2_tvalid ,
	input wire  outport_33_2_tready,
	//output ports STRUCT
	output wire [184-1:0] outport_33_3_tdata ,
	output wire  outport_33_3_tvalid ,
	input wire  outport_33_3_tready,
	//output ports STRUCT
	output wire [112-1:0] outport_33_4_tdata ,
	output wire  outport_33_4_tvalid ,
	input wire  outport_33_4_tready,
	//output ports STRUCT
	output wire [160-1:0] outport_33_5_tdata ,
	output wire  outport_33_5_tvalid ,
	input wire  outport_33_5_tready
);
//
 wire [96-1:0] arg_28_0_tdata;
 wire  arg_28_0_tvalid;
 wire  arg_28_0_tready;

//
 wire [96-1:0] arg_28_1_tdata;
 wire  arg_28_1_tvalid;
 wire  arg_28_1_tready;

//
 wire [96-1:0] arg_28_2_tdata;
 wire  arg_28_2_tvalid;
 wire  arg_28_2_tready;

axis_replication#(
.DATA_WIDTH(96),
.IF_STREAM(0),
.REAPLICA_COUNT(3)
)axis_replication_34(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.s_axis_in_tdata({arg_28_tdata}),
	.s_axis_in_tvalid({arg_28_tvalid}),
	.s_axis_in_tready({arg_28_tready}),
	//
	.m_axis_out_tdata({arg_28_0_tdata,arg_28_1_tdata,arg_28_2_tdata}),
	.m_axis_out_tvalid({arg_28_0_tvalid,arg_28_1_tvalid,arg_28_2_tvalid}),
	.m_axis_out_tready({arg_28_0_tready,arg_28_1_tready,arg_28_2_tready})
);

//const_INT
 wire [32-1:0] const_INT_35_tdata=0;
 wire  const_INT_35_tvalid=1;
 wire  const_INT_35_tready;

//const_INT
 wire [64-1:0] const_INT_36_tdata=0;
 wire  const_INT_36_tvalid=1;
 wire  const_INT_36_tready;

//Table lookup port wire def 
 wire [16-1:0] lookup_p_0_req_index;
 wire  lookup_p_0_req_valid;
 wire  lookup_p_0_req_ready;
 wire  lookup_p_0_value_valid;
 wire  lookup_p_0_value_ready;
 wire [256-1:0] lookup_p_0_value_data;

//Table update port wire def 
 wire [16-1:0] update_p_0_req_index;
 wire  update_p_0_req_index_valid;
 wire  update_p_0_req_index_ready;
 wire [256-1:0] update_p_0_req_data;
 wire  update_p_0_req_data_valid;
 wire  update_p_0_req_data_ready;

cam_arbiter#(
.TABLE_SIZE(16),
.KEY_SIZE(16),
.VALUE_SIZE(256),
.LOOKUP_PORTS(1),
.UPDATE_PORTS(1)
)table_37(
	 .clk(clk), 
	 .rst(rst) ,
	//lookup port 
	.s_lookup_req_index({lookup_p_0_req_index}),
	.s_lookup_req_valid({lookup_p_0_req_valid}),
	.s_lookup_req_ready({lookup_p_0_req_ready}),
	.s_lookup_value_valid({lookup_p_0_value_valid}),
	.s_lookup_value_data({lookup_p_0_value_data}),
	.s_lookup_value_ready({lookup_p_0_value_ready}),
	//update port 
	.s_update_req_index({update_p_0_req_index}),
	.s_update_req_index_valid({update_p_0_req_index_valid}),
	.s_update_req_index_ready({update_p_0_req_index_ready}),
	.s_update_req_data({update_p_0_req_data}),
	.s_update_req_data_valid({update_p_0_req_data_valid}),
	.s_update_req_data_ready({update_p_0_req_data_ready})
);

//Access Struct
 wire [32-1:0] struct_accessed_INT_39_tdata;
 wire  struct_accessed_INT_39_tvalid;
 wire  struct_accessed_INT_39_tready;

struct_access#(
.STRUCT_WIDTH(96),
.ACCESS_OFFSET(0),
.ACCESS_SIZE(32)
)struct_access_38(
	 .clk(clk), 
	 .rst(rst) ,
	//struct input
	.s_struct_axis_tdata({arg_28_0_tdata}),
	.s_struct_axis_tvalid({arg_28_0_tvalid}),
	.s_struct_axis_tready({arg_28_0_tready}),
	//output val
	.m_val_axis_tdata({struct_accessed_INT_39_tdata}),
	.m_val_axis_tvalid({struct_accessed_INT_39_tvalid}),
	.m_val_axis_tready({struct_accessed_INT_39_tready})
);

//bitcast dst
 wire [16-1:0] bitcasted_40_tdata;
 wire  bitcasted_40_tvalid;
 wire  bitcasted_40_tready;

//bitcast dst
 wire [16-1:0] bitcasted_40_0_tdata;
 wire  bitcasted_40_0_tvalid;
 wire  bitcasted_40_0_tready;

//bitcast dst
 wire [16-1:0] bitcasted_40_1_tdata;
 wire  bitcasted_40_1_tvalid;
 wire  bitcasted_40_1_tready;

axis_replication#(
.DATA_WIDTH(16),
.IF_STREAM(0),
.REAPLICA_COUNT(2)
)axis_replication_41(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.s_axis_in_tdata({bitcasted_40_tdata}),
	.s_axis_in_tvalid({bitcasted_40_tvalid}),
	.s_axis_in_tready({bitcasted_40_tready}),
	//
	.m_axis_out_tdata({bitcasted_40_0_tdata,bitcasted_40_1_tdata}),
	.m_axis_out_tvalid({bitcasted_40_0_tvalid,bitcasted_40_1_tvalid}),
	.m_axis_out_tready({bitcasted_40_0_tready,bitcasted_40_1_tready})
);

 assign bitcasted_40_tdata = struct_accessed_INT_39_tdata;
 assign bitcasted_40_tvalid = struct_accessed_INT_39_tvalid;
 assign struct_accessed_INT_39_tready = bitcasted_40_tready;

 assign lookup_p_0_req_index = bitcasted_40_0_tdata;
 assign lookup_p_0_req_valid = bitcasted_40_0_tvalid;
 assign bitcasted_40_0_tready = lookup_p_0_req_ready;

//table lookup resultlookedup_STRUCT_42
 wire [256-1:0] lookedup_STRUCT_42_tdata;
 wire  lookedup_STRUCT_42_tvalid;
 wire  lookedup_STRUCT_42_tready;

//table lookup resultlookedup_STRUCT_42
 wire [256-1:0] lookedup_STRUCT_42_0_tdata;
 wire  lookedup_STRUCT_42_0_tvalid;
 wire  lookedup_STRUCT_42_0_tready;

//table lookup resultlookedup_STRUCT_42
 wire [256-1:0] lookedup_STRUCT_42_1_tdata;
 wire  lookedup_STRUCT_42_1_tvalid;
 wire  lookedup_STRUCT_42_1_tready;

//table lookup resultlookedup_STRUCT_42
 wire [256-1:0] lookedup_STRUCT_42_2_tdata;
 wire  lookedup_STRUCT_42_2_tvalid;
 wire  lookedup_STRUCT_42_2_tready;

//table lookup resultlookedup_STRUCT_42
 wire [256-1:0] lookedup_STRUCT_42_3_tdata;
 wire  lookedup_STRUCT_42_3_tvalid;
 wire  lookedup_STRUCT_42_3_tready;

axis_replication#(
.DATA_WIDTH(256),
.IF_STREAM(0),
.REAPLICA_COUNT(4)
)axis_replication_43(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.s_axis_in_tdata({lookedup_STRUCT_42_tdata}),
	.s_axis_in_tvalid({lookedup_STRUCT_42_tvalid}),
	.s_axis_in_tready({lookedup_STRUCT_42_tready}),
	//
	.m_axis_out_tdata({lookedup_STRUCT_42_0_tdata,lookedup_STRUCT_42_1_tdata,lookedup_STRUCT_42_2_tdata,lookedup_STRUCT_42_3_tdata}),
	.m_axis_out_tvalid({lookedup_STRUCT_42_0_tvalid,lookedup_STRUCT_42_1_tvalid,lookedup_STRUCT_42_2_tvalid,lookedup_STRUCT_42_3_tvalid}),
	.m_axis_out_tready({lookedup_STRUCT_42_0_tready,lookedup_STRUCT_42_1_tready,lookedup_STRUCT_42_2_tready,lookedup_STRUCT_42_3_tready})
);

 assign lookedup_STRUCT_42_tdata = lookup_p_0_value_data;
 assign lookedup_STRUCT_42_tvalid = lookup_p_0_value_valid;
 assign lookup_p_0_value_ready = lookedup_STRUCT_42_tready;

//inited_STRUCT
 wire [96-1:0] inited_STRUCT_44_tdata=0;
 wire  inited_STRUCT_44_tvalid=1;
 wire  inited_STRUCT_44_tready;

//Access Struct
 wire [32-1:0] struct_accessed_INT_46_tdata;
 wire  struct_accessed_INT_46_tvalid;
 wire  struct_accessed_INT_46_tready;

struct_access#(
.STRUCT_WIDTH(256),
.ACCESS_OFFSET(128),
.ACCESS_SIZE(32)
)struct_access_45(
	 .clk(clk), 
	 .rst(rst) ,
	//struct input
	.s_struct_axis_tdata({lookedup_STRUCT_42_0_tdata}),
	.s_struct_axis_tvalid({lookedup_STRUCT_42_0_tvalid}),
	.s_struct_axis_tready({lookedup_STRUCT_42_0_tready}),
	//output val
	.m_val_axis_tdata({struct_accessed_INT_46_tdata}),
	.m_val_axis_tvalid({struct_accessed_INT_46_tvalid}),
	.m_val_axis_tready({struct_accessed_INT_46_tready})
);

//Access Struct
 wire [32-1:0] struct_accessed_INT_48_tdata;
 wire  struct_accessed_INT_48_tvalid;
 wire  struct_accessed_INT_48_tready;

struct_access#(
.STRUCT_WIDTH(96),
.ACCESS_OFFSET(64),
.ACCESS_SIZE(32)
)struct_access_47(
	 .clk(clk), 
	 .rst(rst) ,
	//struct input
	.s_struct_axis_tdata({arg_28_1_tdata}),
	.s_struct_axis_tvalid({arg_28_1_tvalid}),
	.s_struct_axis_tready({arg_28_1_tready}),
	//output val
	.m_val_axis_tdata({struct_accessed_INT_48_tdata}),
	.m_val_axis_tvalid({struct_accessed_INT_48_tvalid}),
	.m_val_axis_tready({struct_accessed_INT_48_tready})
);

//Arithmetic OP Out
 wire [32-1:0] SUB_49_out_INT_50_tdata = 0;
 wire  SUB_49_out_INT_50_tvalid;
 wire  SUB_49_out_INT_50_tready;

//Arithmetic OP Out
 wire [32-1:0] SUB_49_out_INT_50_0_tdata;
 wire  SUB_49_out_INT_50_0_tvalid;
 wire  SUB_49_out_INT_50_0_tready;

//Arithmetic OP Out
 wire [32-1:0] SUB_49_out_INT_50_1_tdata;
 wire  SUB_49_out_INT_50_1_tvalid;
 wire  SUB_49_out_INT_50_1_tready;

//Arithmetic OP Out
 wire [32-1:0] SUB_49_out_INT_50_2_tdata;
 wire  SUB_49_out_INT_50_2_tvalid;
 wire  SUB_49_out_INT_50_2_tready;

axis_replication#(
.DATA_WIDTH(32),
.IF_STREAM(0),
.REAPLICA_COUNT(3)
)axis_replication_51(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.s_axis_in_tdata({SUB_49_out_INT_50_tdata}),
	.s_axis_in_tvalid({SUB_49_out_INT_50_tvalid}),
	.s_axis_in_tready({SUB_49_out_INT_50_tready}),
	//
	.m_axis_out_tdata({SUB_49_out_INT_50_0_tdata,SUB_49_out_INT_50_1_tdata,SUB_49_out_INT_50_2_tdata}),
	.m_axis_out_tvalid({SUB_49_out_INT_50_0_tvalid,SUB_49_out_INT_50_1_tvalid,SUB_49_out_INT_50_2_tvalid}),
	.m_axis_out_tready({SUB_49_out_INT_50_0_tready,SUB_49_out_INT_50_1_tready,SUB_49_out_INT_50_2_tready})
);

ALU#(
.LVAL_SIZE(32),
.RVAL_SIZE(32),
.RESULT_SIZE(32),
.OPID(0)
)SUB_49(
	 .clk(clk), 
	 .rst(rst) ,
	//lval input
	.s_lval_axis_tdata({struct_accessed_INT_46_tdata}),
	.s_lval_axis_tvalid({struct_accessed_INT_46_tvalid}),
	.s_lval_axis_tready({struct_accessed_INT_46_tready}),
	//rval input
	.s_rval_axis_tdata({struct_accessed_INT_48_tdata}),
	.s_rval_axis_tvalid({struct_accessed_INT_48_tvalid}),
	.s_rval_axis_tready({struct_accessed_INT_48_tready}),
	//output val
	.m_val_axis_tdata({}),
	.m_val_axis_tvalid({SUB_49_out_INT_50_tvalid}),
	.m_val_axis_tready({SUB_49_out_INT_50_tready})
);

//Access Struct
 wire [32-1:0] struct_accessed_INT_53_tdata;
 wire  struct_accessed_INT_53_tvalid;
 wire  struct_accessed_INT_53_tready;

//Access Struct
 wire [32-1:0] struct_accessed_INT_53_0_tdata;
 wire  struct_accessed_INT_53_0_tvalid;
 wire  struct_accessed_INT_53_0_tready;

//Access Struct
 wire [32-1:0] struct_accessed_INT_53_1_tdata;
 wire  struct_accessed_INT_53_1_tvalid;
 wire  struct_accessed_INT_53_1_tready;

//Access Struct
 wire [32-1:0] struct_accessed_INT_53_2_tdata;
 wire  struct_accessed_INT_53_2_tvalid;
 wire  struct_accessed_INT_53_2_tready;

axis_replication#(
.DATA_WIDTH(32),
.IF_STREAM(0),
.REAPLICA_COUNT(3)
)axis_replication_54(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.s_axis_in_tdata({struct_accessed_INT_53_tdata}),
	.s_axis_in_tvalid({struct_accessed_INT_53_tvalid}),
	.s_axis_in_tready({struct_accessed_INT_53_tready}),
	//
	.m_axis_out_tdata({struct_accessed_INT_53_0_tdata,struct_accessed_INT_53_1_tdata,struct_accessed_INT_53_2_tdata}),
	.m_axis_out_tvalid({struct_accessed_INT_53_0_tvalid,struct_accessed_INT_53_1_tvalid,struct_accessed_INT_53_2_tvalid}),
	.m_axis_out_tready({struct_accessed_INT_53_0_tready,struct_accessed_INT_53_1_tready,struct_accessed_INT_53_2_tready})
);

struct_access#(
.STRUCT_WIDTH(96),
.ACCESS_OFFSET(32),
.ACCESS_SIZE(32)
)struct_access_52(
	 .clk(clk), 
	 .rst(rst) ,
	//struct input
	.s_struct_axis_tdata({arg_28_2_tdata}),
	.s_struct_axis_tvalid({arg_28_2_tvalid}),
	.s_struct_axis_tready({arg_28_2_tready}),
	//output val
	.m_val_axis_tdata({struct_accessed_INT_53_tdata}),
	.m_val_axis_tvalid({struct_accessed_INT_53_tvalid}),
	.m_val_axis_tready({struct_accessed_INT_53_tready})
);

//Arithmetic OP Out
 wire [32-1:0] SUB_55_out_INT_56_tdata;
 wire  SUB_55_out_INT_56_tvalid;
 wire  SUB_55_out_INT_56_tready;

//Arithmetic OP Out
 wire [32-1:0] SUB_55_out_INT_56_0_tdata;
 wire  SUB_55_out_INT_56_0_tvalid;
 wire  SUB_55_out_INT_56_0_tready;

//Arithmetic OP Out
 wire [32-1:0] SUB_55_out_INT_56_1_tdata;
 wire  SUB_55_out_INT_56_1_tvalid;
 wire  SUB_55_out_INT_56_1_tready;

axis_replication#(
.DATA_WIDTH(32),
.IF_STREAM(0),
.REAPLICA_COUNT(2)
)axis_replication_57(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.s_axis_in_tdata({SUB_55_out_INT_56_tdata}),
	.s_axis_in_tvalid({SUB_55_out_INT_56_tvalid}),
	.s_axis_in_tready({SUB_55_out_INT_56_tready}),
	//
	.m_axis_out_tdata({SUB_55_out_INT_56_0_tdata,SUB_55_out_INT_56_1_tdata}),
	.m_axis_out_tvalid({SUB_55_out_INT_56_0_tvalid,SUB_55_out_INT_56_1_tvalid}),
	.m_axis_out_tready({SUB_55_out_INT_56_0_tready,SUB_55_out_INT_56_1_tready})
);

ALU#(
.LVAL_SIZE(32),
.RVAL_SIZE(32),
.RESULT_SIZE(32),
.OPID(0)
)SUB_55(
	 .clk(clk), 
	 .rst(rst) ,
	//lval input
	.s_lval_axis_tdata({struct_accessed_INT_53_0_tdata}),
	.s_lval_axis_tvalid({struct_accessed_INT_53_0_tvalid}),
	.s_lval_axis_tready({struct_accessed_INT_53_0_tready}),
	//rval input
	.s_rval_axis_tdata({SUB_49_out_INT_50_0_tdata}),
	.s_rval_axis_tvalid({SUB_49_out_INT_50_0_tvalid}),
	.s_rval_axis_tready({SUB_49_out_INT_50_0_tready}),
	//output val
	.m_val_axis_tdata({SUB_55_out_INT_56_tdata}),
	.m_val_axis_tvalid({SUB_55_out_INT_56_tvalid}),
	.m_val_axis_tready({SUB_55_out_INT_56_tready})
);

//Access Struct
 wire [32-1:0] struct_accessed_INT_59_tdata;
 wire  struct_accessed_INT_59_tvalid;
 wire  struct_accessed_INT_59_tready;

//Access Struct
 wire [32-1:0] struct_accessed_INT_59_0_tdata;
 wire  struct_accessed_INT_59_0_tvalid;
 wire  struct_accessed_INT_59_0_tready;

//Access Struct
 wire [32-1:0] struct_accessed_INT_59_1_tdata;
 wire  struct_accessed_INT_59_1_tvalid;
 wire  struct_accessed_INT_59_1_tready;

//Access Struct
 wire [32-1:0] struct_accessed_INT_59_2_tdata;
 wire  struct_accessed_INT_59_2_tvalid;
 wire  struct_accessed_INT_59_2_tready;

axis_replication#(
.DATA_WIDTH(32),
.IF_STREAM(0),
.REAPLICA_COUNT(3)
)axis_replication_60(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.s_axis_in_tdata({struct_accessed_INT_59_tdata}),
	.s_axis_in_tvalid({struct_accessed_INT_59_tvalid}),
	.s_axis_in_tready({struct_accessed_INT_59_tready}),
	//
	.m_axis_out_tdata({struct_accessed_INT_59_0_tdata,struct_accessed_INT_59_1_tdata,struct_accessed_INT_59_2_tdata}),
	.m_axis_out_tvalid({struct_accessed_INT_59_0_tvalid,struct_accessed_INT_59_1_tvalid,struct_accessed_INT_59_2_tvalid}),
	.m_axis_out_tready({struct_accessed_INT_59_0_tready,struct_accessed_INT_59_1_tready,struct_accessed_INT_59_2_tready})
);

struct_access#(
.STRUCT_WIDTH(256),
.ACCESS_OFFSET(96),
.ACCESS_SIZE(32)
)struct_access_58(
	 .clk(clk), 
	 .rst(rst) ,
	//struct input
	.s_struct_axis_tdata({lookedup_STRUCT_42_1_tdata}),
	.s_struct_axis_tvalid({lookedup_STRUCT_42_1_tvalid}),
	.s_struct_axis_tready({lookedup_STRUCT_42_1_tready}),
	//output val
	.m_val_axis_tdata({struct_accessed_INT_59_tdata}),
	.m_val_axis_tvalid({struct_accessed_INT_59_tvalid}),
	.m_val_axis_tready({struct_accessed_INT_59_tready})
);

//Arithmetic OP Out
 wire [1-1:0] LT_61_out_INT_62_tdata;
 wire  LT_61_out_INT_62_tvalid;
 wire  LT_61_out_INT_62_tready;

ALU#(
.LVAL_SIZE(32),
.RVAL_SIZE(32),
.RESULT_SIZE(1),
.OPID(3)
)LT_61(
	 .clk(clk), 
	 .rst(rst) ,
	//lval input
	.s_lval_axis_tdata({SUB_55_out_INT_56_0_tdata}),
	.s_lval_axis_tvalid({SUB_55_out_INT_56_0_tvalid}),
	.s_lval_axis_tready({SUB_55_out_INT_56_0_tready}),
	//rval input
	.s_rval_axis_tdata({struct_accessed_INT_59_0_tdata}),
	.s_rval_axis_tvalid({struct_accessed_INT_59_0_tvalid}),
	.s_rval_axis_tready({struct_accessed_INT_59_0_tready}),
	//output val
	.m_val_axis_tdata({LT_61_out_INT_62_tdata}),
	.m_val_axis_tvalid({LT_61_out_INT_62_tvalid}),
	.m_val_axis_tready({LT_61_out_INT_62_tready})
);

//Arithmetic OP Out
 wire [32-1:0] SUB_63_out_INT_64_tdata;
 wire  SUB_63_out_INT_64_tvalid;
 wire  SUB_63_out_INT_64_tready;

ALU#(
.LVAL_SIZE(32),
.RVAL_SIZE(32),
.RESULT_SIZE(32),
.OPID(0)
)SUB_63(
	 .clk(clk), 
	 .rst(rst) ,
	//lval input
	.s_lval_axis_tdata({SUB_55_out_INT_56_1_tdata}),
	.s_lval_axis_tvalid({SUB_55_out_INT_56_1_tvalid}),
	.s_lval_axis_tready({SUB_55_out_INT_56_1_tready}),
	//rval input
	.s_rval_axis_tdata({struct_accessed_INT_59_1_tdata}),
	.s_rval_axis_tvalid({struct_accessed_INT_59_1_tvalid}),
	.s_rval_axis_tready({struct_accessed_INT_59_1_tready}),
	//output val
	.m_val_axis_tdata({SUB_63_out_INT_64_tdata}),
	.m_val_axis_tvalid({SUB_63_out_INT_64_tvalid}),
	.m_val_axis_tready({SUB_63_out_INT_64_tready})
);

//Arithmetic OP Out
 wire [1-1:0] LE_65_out_INT_66_tdata;
 wire  LE_65_out_INT_66_tvalid;
 wire  LE_65_out_INT_66_tready;

//Arithmetic OP Out
 wire [1-1:0] LE_65_out_INT_66_0_tdata;
 wire  LE_65_out_INT_66_0_tvalid;
 wire  LE_65_out_INT_66_0_tready;

//Arithmetic OP Out
 wire [1-1:0] LE_65_out_INT_66_1_tdata;
 wire  LE_65_out_INT_66_1_tvalid;
 wire  LE_65_out_INT_66_1_tready;

axis_replication#(
.DATA_WIDTH(1),
.IF_STREAM(0),
.REAPLICA_COUNT(2)
)axis_replication_67(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.s_axis_in_tdata({LE_65_out_INT_66_tdata}),
	.s_axis_in_tvalid({LE_65_out_INT_66_tvalid}),
	.s_axis_in_tready({LE_65_out_INT_66_tready}),
	//
	.m_axis_out_tdata({LE_65_out_INT_66_0_tdata,LE_65_out_INT_66_1_tdata}),
	.m_axis_out_tvalid({LE_65_out_INT_66_0_tvalid,LE_65_out_INT_66_1_tvalid}),
	.m_axis_out_tready({LE_65_out_INT_66_0_tready,LE_65_out_INT_66_1_tready})
);

ALU#(
.LVAL_SIZE(32),
.RVAL_SIZE(32),
.RESULT_SIZE(1),
.OPID(6)
)LE_65(
	 .clk(clk), 
	 .rst(rst) ,
	//lval input
	.s_lval_axis_tdata({SUB_49_out_INT_50_1_tdata}),
	.s_lval_axis_tvalid({SUB_49_out_INT_50_1_tvalid}),
	.s_lval_axis_tready({SUB_49_out_INT_50_1_tready}),
	//rval input
	.s_rval_axis_tdata({struct_accessed_INT_53_1_tdata}),
	.s_rval_axis_tvalid({struct_accessed_INT_53_1_tvalid}),
	.s_rval_axis_tready({struct_accessed_INT_53_1_tready}),
	//output val
	.m_val_axis_tdata({LE_65_out_INT_66_tdata}),
	.m_val_axis_tvalid({LE_65_out_INT_66_tvalid}),
	.m_val_axis_tready({LE_65_out_INT_66_tready})
);

//
 wire [32-1:0] select_result_68_tdata;
 wire  select_result_68_tvalid;
 wire  select_result_68_tready;

select#(
.VAL_WIDTH(32),
.COND_WIDTH(1)
)select_69(
	 .clk(clk), 
	 .rst(rst) ,
	//select condition
	.s_cond_axis_tdata({LT_61_out_INT_62_tdata}),
	.s_cond_axis_tvalid({LT_61_out_INT_62_tvalid}),
	.s_cond_axis_tready({LT_61_out_INT_62_tready}),
	//select true val
	.s_true_val_axis_tdata({const_INT_35_tdata}),
	.s_true_val_axis_tvalid({const_INT_35_tvalid}),
	.s_true_val_axis_tready({const_INT_35_tready}),
	//select false val
	.s_false_val_axis_tdata({SUB_63_out_INT_64_tdata}),
	.s_false_val_axis_tvalid({SUB_63_out_INT_64_tvalid}),
	.s_false_val_axis_tready({SUB_63_out_INT_64_tready}),
	//select result
	.m_val_axis_tdata({select_result_68_tdata}),
	.m_val_axis_tvalid({select_result_68_tvalid}),
	.m_val_axis_tready({select_result_68_tready})
);

//Arithmetic OP Out
 wire [32-1:0] ADD_70_out_INT_71_tdata;
 wire  ADD_70_out_INT_71_tvalid;
 wire  ADD_70_out_INT_71_tready;

ALU#(
.LVAL_SIZE(32),
.RVAL_SIZE(32),
.RESULT_SIZE(32),
.OPID(1)
)ADD_70(
	 .clk(clk), 
	 .rst(rst) ,
	//lval input
	.s_lval_axis_tdata({SUB_49_out_INT_50_2_tdata}),
	.s_lval_axis_tvalid({SUB_49_out_INT_50_2_tvalid}),
	.s_lval_axis_tready({SUB_49_out_INT_50_2_tready}),
	//rval input
	.s_rval_axis_tdata({select_result_68_tdata}),
	.s_rval_axis_tvalid({select_result_68_tvalid}),
	.s_rval_axis_tready({select_result_68_tready}),
	//output val
	.m_val_axis_tdata({ADD_70_out_INT_71_tdata}),
	.m_val_axis_tvalid({ADD_70_out_INT_71_tvalid}),
	.m_val_axis_tready({ADD_70_out_INT_71_tready})
);

//Arithmetic OP Out
 wire [32-1:0] SUB_72_out_INT_73_tdata;
 wire  SUB_72_out_INT_73_tvalid;
 wire  SUB_72_out_INT_73_tready;

//Arithmetic OP Out
 wire [32-1:0] SUB_72_out_INT_73_0_tdata;
 wire  SUB_72_out_INT_73_0_tvalid;
 wire  SUB_72_out_INT_73_0_tready;

//Arithmetic OP Out
 wire [32-1:0] SUB_72_out_INT_73_1_tdata;
 wire  SUB_72_out_INT_73_1_tvalid;
 wire  SUB_72_out_INT_73_1_tready;

//Arithmetic OP Out
 wire [32-1:0] SUB_72_out_INT_73_2_tdata;
 wire  SUB_72_out_INT_73_2_tvalid;
 wire  SUB_72_out_INT_73_2_tready;

//Arithmetic OP Out
 wire [32-1:0] SUB_72_out_INT_73_3_tdata;
 wire  SUB_72_out_INT_73_3_tvalid;
 wire  SUB_72_out_INT_73_3_tready;

axis_replication#(
.DATA_WIDTH(32),
.IF_STREAM(0),
.REAPLICA_COUNT(4)
)axis_replication_74(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.s_axis_in_tdata({SUB_72_out_INT_73_tdata}),
	.s_axis_in_tvalid({SUB_72_out_INT_73_tvalid}),
	.s_axis_in_tready({SUB_72_out_INT_73_tready}),
	//
	.m_axis_out_tdata({SUB_72_out_INT_73_0_tdata,SUB_72_out_INT_73_1_tdata,SUB_72_out_INT_73_2_tdata,SUB_72_out_INT_73_3_tdata}),
	.m_axis_out_tvalid({SUB_72_out_INT_73_0_tvalid,SUB_72_out_INT_73_1_tvalid,SUB_72_out_INT_73_2_tvalid,SUB_72_out_INT_73_3_tvalid}),
	.m_axis_out_tready({SUB_72_out_INT_73_0_tready,SUB_72_out_INT_73_1_tready,SUB_72_out_INT_73_2_tready,SUB_72_out_INT_73_3_tready})
);

ALU#(
.LVAL_SIZE(32),
.RVAL_SIZE(32),
.RESULT_SIZE(32),
.OPID(0)
)SUB_72(
	 .clk(clk), 
	 .rst(rst) ,
	//lval input
	.s_lval_axis_tdata({struct_accessed_INT_53_2_tdata}),
	.s_lval_axis_tvalid({struct_accessed_INT_53_2_tvalid}),
	.s_lval_axis_tready({struct_accessed_INT_53_2_tready}),
	//rval input
	.s_rval_axis_tdata({ADD_70_out_INT_71_tdata}),
	.s_rval_axis_tvalid({ADD_70_out_INT_71_tvalid}),
	.s_rval_axis_tready({ADD_70_out_INT_71_tready}),
	//output val
	.m_val_axis_tdata({SUB_72_out_INT_73_tdata}),
	.m_val_axis_tvalid({SUB_72_out_INT_73_tvalid}),
	.m_val_axis_tready({SUB_72_out_INT_73_tready})
);

//Arithmetic OP Out
 wire [1-1:0] GT_75_out_INT_76_tdata;
 wire  GT_75_out_INT_76_tvalid;
 wire  GT_75_out_INT_76_tready;

ALU#(
.LVAL_SIZE(32),
.RVAL_SIZE(64),
.RESULT_SIZE(1),
.OPID(4)
)GT_75(
	 .clk(clk), 
	 .rst(rst) ,
	//lval input
	.s_lval_axis_tdata({SUB_72_out_INT_73_0_tdata}),
	.s_lval_axis_tvalid({SUB_72_out_INT_73_0_tvalid}),
	.s_lval_axis_tready({SUB_72_out_INT_73_0_tready}),
	//rval input
	.s_rval_axis_tdata({const_INT_36_tdata}),
	.s_rval_axis_tvalid({const_INT_36_tvalid}),
	.s_rval_axis_tready({const_INT_36_tready}),
	//output val
	.m_val_axis_tdata({GT_75_out_INT_76_tdata}),
	.m_val_axis_tvalid({GT_75_out_INT_76_tvalid}),
	.m_val_axis_tready({GT_75_out_INT_76_tready})
);

//Arithmetic OP Out
 wire [32-1:0] SUB_77_out_INT_78_tdata;
 wire  SUB_77_out_INT_78_tvalid;
 wire  SUB_77_out_INT_78_tready;

ALU#(
.LVAL_SIZE(32),
.RVAL_SIZE(32),
.RESULT_SIZE(32),
.OPID(0)
)SUB_77(
	 .clk(clk), 
	 .rst(rst) ,
	//lval input
	.s_lval_axis_tdata({struct_accessed_INT_59_2_tdata}),
	.s_lval_axis_tvalid({struct_accessed_INT_59_2_tvalid}),
	.s_lval_axis_tready({struct_accessed_INT_59_2_tready}),
	//rval input
	.s_rval_axis_tdata({SUB_72_out_INT_73_1_tdata}),
	.s_rval_axis_tvalid({SUB_72_out_INT_73_1_tvalid}),
	.s_rval_axis_tready({SUB_72_out_INT_73_1_tready}),
	//output val
	.m_val_axis_tdata({SUB_77_out_INT_78_tdata}),
	.m_val_axis_tvalid({SUB_77_out_INT_78_tvalid}),
	.m_val_axis_tready({SUB_77_out_INT_78_tready})
);

//struct_assign_79 output struct
 wire [256-1:0] structvar_80_tdata;
 wire  structvar_80_tvalid;
 wire  structvar_80_tready;

//struct_assign_79 output struct
 wire [256-1:0] structvar_80_0_tdata;
 wire  structvar_80_0_tvalid;
 wire  structvar_80_0_tready;

//struct_assign_79 output struct
 wire [256-1:0] structvar_80_1_tdata;
 wire  structvar_80_1_tvalid;
 wire  structvar_80_1_tready;

axis_replication#(
.DATA_WIDTH(256),
.IF_STREAM(0),
.REAPLICA_COUNT(2)
)axis_replication_81(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.s_axis_in_tdata({structvar_80_tdata}),
	.s_axis_in_tvalid({structvar_80_tvalid}),
	.s_axis_in_tready({structvar_80_tready}),
	//
	.m_axis_out_tdata({structvar_80_0_tdata,structvar_80_1_tdata}),
	.m_axis_out_tvalid({structvar_80_0_tvalid,structvar_80_1_tvalid}),
	.m_axis_out_tready({structvar_80_0_tready,structvar_80_1_tready})
);

struct_assign#(
.STRUCT_WIDTH(256),
.ASSIGN_OFFSET(96),
.ASSIGN_SIZE(32)
)struct_assign_79(
	 .clk(clk), 
	 .rst(rst) ,
	//input struct
	.s_struct_axis_tdata({lookedup_STRUCT_42_2_tdata}),
	.s_struct_axis_tvalid({lookedup_STRUCT_42_2_tvalid}),
	.s_struct_axis_tready({lookedup_STRUCT_42_2_tready}),
	//input val
	.s_assignv_axis_tdata({SUB_77_out_INT_78_tdata}),
	.s_assignv_axis_tvalid({SUB_77_out_INT_78_tvalid}),
	.s_assignv_axis_tready({SUB_77_out_INT_78_tready}),
	//output struct
	.m_struct_axis_tdata({structvar_80_tdata}),
	.m_struct_axis_tvalid({structvar_80_tvalid}),
	.m_struct_axis_tready({structvar_80_tready})
);

//Access Struct
 wire [32-1:0] struct_accessed_INT_83_tdata;
 wire  struct_accessed_INT_83_tvalid;
 wire  struct_accessed_INT_83_tready;

struct_access#(
.STRUCT_WIDTH(256),
.ACCESS_OFFSET(128),
.ACCESS_SIZE(32)
)struct_access_82(
	 .clk(clk), 
	 .rst(rst) ,
	//struct input
	.s_struct_axis_tdata({structvar_80_0_tdata}),
	.s_struct_axis_tvalid({structvar_80_0_tvalid}),
	.s_struct_axis_tready({structvar_80_0_tready}),
	//output val
	.m_val_axis_tdata({struct_accessed_INT_83_tdata}),
	.m_val_axis_tvalid({struct_accessed_INT_83_tvalid}),
	.m_val_axis_tready({struct_accessed_INT_83_tready})
);

//Arithmetic OP Out
 wire [32-1:0] ADD_84_out_INT_85_tdata;
 wire  ADD_84_out_INT_85_tvalid;
 wire  ADD_84_out_INT_85_tready;

ALU#(
.LVAL_SIZE(32),
.RVAL_SIZE(32),
.RESULT_SIZE(32),
.OPID(1)
)ADD_84(
	 .clk(clk), 
	 .rst(rst) ,
	//lval input
	.s_lval_axis_tdata({struct_accessed_INT_83_tdata}),
	.s_lval_axis_tvalid({struct_accessed_INT_83_tvalid}),
	.s_lval_axis_tready({struct_accessed_INT_83_tready}),
	//rval input
	.s_rval_axis_tdata({SUB_72_out_INT_73_2_tdata}),
	.s_rval_axis_tvalid({SUB_72_out_INT_73_2_tvalid}),
	.s_rval_axis_tready({SUB_72_out_INT_73_2_tready}),
	//output val
	.m_val_axis_tdata({ADD_84_out_INT_85_tdata}),
	.m_val_axis_tvalid({ADD_84_out_INT_85_tvalid}),
	.m_val_axis_tready({ADD_84_out_INT_85_tready})
);

//struct_assign_86 output struct
 wire [256-1:0] structvar_87_tdata;
 wire  structvar_87_tvalid;
 wire  structvar_87_tready;

//struct_assign_86 output struct
 wire [256-1:0] structvar_87_0_tdata;
 wire  structvar_87_0_tvalid;
 wire  structvar_87_0_tready;

//struct_assign_86 output struct
 wire [256-1:0] structvar_87_1_tdata;
 wire  structvar_87_1_tvalid;
 wire  structvar_87_1_tready;

axis_replication#(
.DATA_WIDTH(256),
.IF_STREAM(0),
.REAPLICA_COUNT(2)
)axis_replication_88(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.s_axis_in_tdata({structvar_87_tdata}),
	.s_axis_in_tvalid({structvar_87_tvalid}),
	.s_axis_in_tready({structvar_87_tready}),
	//
	.m_axis_out_tdata({structvar_87_0_tdata,structvar_87_1_tdata}),
	.m_axis_out_tvalid({structvar_87_0_tvalid,structvar_87_1_tvalid}),
	.m_axis_out_tready({structvar_87_0_tready,structvar_87_1_tready})
);

struct_assign#(
.STRUCT_WIDTH(256),
.ASSIGN_OFFSET(128),
.ASSIGN_SIZE(32)
)struct_assign_86(
	 .clk(clk), 
	 .rst(rst) ,
	//input struct
	.s_struct_axis_tdata({structvar_80_1_tdata}),
	.s_struct_axis_tvalid({structvar_80_1_tvalid}),
	.s_struct_axis_tready({structvar_80_1_tready}),
	//input val
	.s_assignv_axis_tdata({ADD_84_out_INT_85_tdata}),
	.s_assignv_axis_tvalid({ADD_84_out_INT_85_tvalid}),
	.s_assignv_axis_tready({ADD_84_out_INT_85_tready}),
	//output struct
	.m_struct_axis_tdata({structvar_87_tdata}),
	.m_struct_axis_tvalid({structvar_87_tvalid}),
	.m_struct_axis_tready({structvar_87_tready})
);

//Access Struct
 wire [32-1:0] struct_accessed_INT_90_tdata;
 wire  struct_accessed_INT_90_tvalid;
 wire  struct_accessed_INT_90_tready;

struct_access#(
.STRUCT_WIDTH(256),
.ACCESS_OFFSET(160),
.ACCESS_SIZE(32)
)struct_access_89(
	 .clk(clk), 
	 .rst(rst) ,
	//struct input
	.s_struct_axis_tdata({structvar_87_0_tdata}),
	.s_struct_axis_tvalid({structvar_87_0_tvalid}),
	.s_struct_axis_tready({structvar_87_0_tready}),
	//output val
	.m_val_axis_tdata({struct_accessed_INT_90_tdata}),
	.m_val_axis_tvalid({struct_accessed_INT_90_tvalid}),
	.m_val_axis_tready({struct_accessed_INT_90_tready})
);

//Arithmetic OP Out
 wire [32-1:0] ADD_91_out_INT_92_tdata;
 wire  ADD_91_out_INT_92_tvalid;
 wire  ADD_91_out_INT_92_tready;

ALU#(
.LVAL_SIZE(32),
.RVAL_SIZE(32),
.RESULT_SIZE(32),
.OPID(1)
)ADD_91(
	 .clk(clk), 
	 .rst(rst) ,
	//lval input
	.s_lval_axis_tdata({struct_accessed_INT_90_tdata}),
	.s_lval_axis_tvalid({struct_accessed_INT_90_tvalid}),
	.s_lval_axis_tready({struct_accessed_INT_90_tready}),
	//rval input
	.s_rval_axis_tdata({SUB_72_out_INT_73_3_tdata}),
	.s_rval_axis_tvalid({SUB_72_out_INT_73_3_tvalid}),
	.s_rval_axis_tready({SUB_72_out_INT_73_3_tready}),
	//output val
	.m_val_axis_tdata({ADD_91_out_INT_92_tdata}),
	.m_val_axis_tvalid({ADD_91_out_INT_92_tvalid}),
	.m_val_axis_tready({ADD_91_out_INT_92_tready})
);

//struct_assign_93 output struct
 wire [256-1:0] structvar_94_tdata;
 wire  structvar_94_tvalid;
 wire  structvar_94_tready;

struct_assign#(
.STRUCT_WIDTH(256),
.ASSIGN_OFFSET(160),
.ASSIGN_SIZE(32)
)struct_assign_93(
	 .clk(clk), 
	 .rst(rst) ,
	//input struct
	.s_struct_axis_tdata({structvar_87_1_tdata}),
	.s_struct_axis_tvalid({structvar_87_1_tvalid}),
	.s_struct_axis_tready({structvar_87_1_tready}),
	//input val
	.s_assignv_axis_tdata({ADD_91_out_INT_92_tdata}),
	.s_assignv_axis_tvalid({ADD_91_out_INT_92_tvalid}),
	.s_assignv_axis_tready({ADD_91_out_INT_92_tready}),
	//output struct
	.m_struct_axis_tdata({structvar_94_tdata}),
	.m_struct_axis_tvalid({structvar_94_tvalid}),
	.m_struct_axis_tready({structvar_94_tready})
);

//
 wire [256-1:0] select_result_95_tdata;
 wire  select_result_95_tvalid;
 wire  select_result_95_tready;

//
 wire [256-1:0] select_result_95_0_tdata;
 wire  select_result_95_0_tvalid;
 wire  select_result_95_0_tready;

//
 wire [256-1:0] select_result_95_1_tdata;
 wire  select_result_95_1_tvalid;
 wire  select_result_95_1_tready;

//
 wire [256-1:0] select_result_95_2_tdata;
 wire  select_result_95_2_tvalid;
 wire  select_result_95_2_tready;

//
 wire [256-1:0] select_result_95_3_tdata;
 wire  select_result_95_3_tvalid;
 wire  select_result_95_3_tready;

axis_replication#(
.DATA_WIDTH(256),
.IF_STREAM(0),
.REAPLICA_COUNT(4)
)axis_replication_96(
	 .clk(clk), 
	 .rst(rst) ,
	//
	.s_axis_in_tdata({select_result_95_tdata}),
	.s_axis_in_tvalid({select_result_95_tvalid}),
	.s_axis_in_tready({select_result_95_tready}),
	//
	.m_axis_out_tdata({select_result_95_0_tdata,select_result_95_1_tdata,select_result_95_2_tdata,select_result_95_3_tdata}),
	.m_axis_out_tvalid({select_result_95_0_tvalid,select_result_95_1_tvalid,select_result_95_2_tvalid,select_result_95_3_tvalid}),
	.m_axis_out_tready({select_result_95_0_tready,select_result_95_1_tready,select_result_95_2_tready,select_result_95_3_tready})
);

select#(
.VAL_WIDTH(256),
.COND_WIDTH(1)
)select_97(
	 .clk(clk), 
	 .rst(rst) ,
	//select condition
	.s_cond_axis_tdata({GT_75_out_INT_76_tdata}),
	.s_cond_axis_tvalid({GT_75_out_INT_76_tvalid}),
	.s_cond_axis_tready({GT_75_out_INT_76_tready}),
	//select true val
	.s_true_val_axis_tdata({structvar_94_tdata}),
	.s_true_val_axis_tvalid({structvar_94_tvalid}),
	.s_true_val_axis_tready({structvar_94_tready}),
	//select false val
	.s_false_val_axis_tdata({lookedup_STRUCT_42_3_tdata}),
	.s_false_val_axis_tvalid({lookedup_STRUCT_42_3_tvalid}),
	.s_false_val_axis_tready({lookedup_STRUCT_42_3_tready}),
	//select result
	.m_val_axis_tdata({select_result_95_tdata}),
	.m_val_axis_tvalid({select_result_95_tvalid}),
	.m_val_axis_tready({select_result_95_tready})
);

//replicated guard condition
 wire [1-1:0] replicated_guard_cond_98_tdata;
 wire  replicated_guard_cond_98_tvalid;
 wire  replicated_guard_cond_98_tready;

//replicated guard condition
 wire [1-1:0] replicated_guard_cond_99_tdata;
 wire  replicated_guard_cond_99_tvalid;
 wire  replicated_guard_cond_99_tready;

guard_pred#(
.COND_WIDTH(1),
.REPLICATED_OUT_NUM(2),
.GROUND_TRUTH(1)
)guard_pred_100(
	 .clk(clk), 
	 .rst(rst) ,
	//guard condition
	.s_guard_cond_tdata({LE_65_out_INT_66_0_tdata}),
	.s_guard_cond_tvalid({LE_65_out_INT_66_0_tvalid}),
	.s_guard_cond_tready({LE_65_out_INT_66_0_tready}),
	//replicated guard condition
	.m_guard_cond_tdata({replicated_guard_cond_98_tdata,replicated_guard_cond_99_tdata}),
	.m_guard_cond_tvalid({replicated_guard_cond_98_tvalid,replicated_guard_cond_99_tvalid}),
	.m_guard_cond_tready({replicated_guard_cond_98_tready,replicated_guard_cond_99_tready})
);

//-- guarded
 wire [16-1:0] bitcasted_40_1_guarded_tdata;
 wire  bitcasted_40_1_guarded_tvalid;
 wire  bitcasted_40_1_guarded_tready;

guard#(
.DATA_WIDTH(16),
.IF_STREAM(0)
)guard_101(
	 .clk(clk), 
	 .rst(rst) ,
	//input val
	.s_guard_axis_tdata({bitcasted_40_1_tdata}),
	.s_guard_axis_tvalid({bitcasted_40_1_tvalid}),
	.s_guard_axis_tready({bitcasted_40_1_tready}),
	//output val
	.m_guard_axis_tdata({bitcasted_40_1_guarded_tdata}),
	.m_guard_axis_tvalid({bitcasted_40_1_guarded_tvalid}),
	.m_guard_axis_tready({bitcasted_40_1_guarded_tready}),
	//guard condition
	.s_guard_cond_tdata({replicated_guard_cond_98_tdata}),
	.s_guard_cond_tvalid({replicated_guard_cond_98_tvalid}),
	.s_guard_cond_tready({replicated_guard_cond_98_tready})
);

//-- guarded
 wire [256-1:0] select_result_95_0_guarded_tdata;
 wire  select_result_95_0_guarded_tvalid;
 wire  select_result_95_0_guarded_tready;

guard#(
.DATA_WIDTH(256),
.IF_STREAM(0)
)guard_102(
	 .clk(clk), 
	 .rst(rst) ,
	//input val
	.s_guard_axis_tdata({select_result_95_0_tdata}),
	.s_guard_axis_tvalid({select_result_95_0_tvalid}),
	.s_guard_axis_tready({select_result_95_0_tready}),
	//output val
	.m_guard_axis_tdata({select_result_95_0_guarded_tdata}),
	.m_guard_axis_tvalid({select_result_95_0_guarded_tvalid}),
	.m_guard_axis_tready({select_result_95_0_guarded_tready}),
	//guard condition
	.s_guard_cond_tdata({replicated_guard_cond_99_tdata}),
	.s_guard_cond_tvalid({replicated_guard_cond_99_tvalid}),
	.s_guard_cond_tready({replicated_guard_cond_99_tready})
);

 assign update_p_0_req_index = bitcasted_40_1_guarded_tdata;
 assign update_p_0_req_index_valid = bitcasted_40_1_guarded_tvalid;
 assign bitcasted_40_1_guarded_tready = update_p_0_req_index_ready;

 assign update_p_0_req_data = select_result_95_0_guarded_tdata;
 assign update_p_0_req_data_valid = select_result_95_0_guarded_tvalid;
 assign select_result_95_0_guarded_tready = update_p_0_req_data_ready;

//Access Struct
 wire [32-1:0] struct_accessed_INT_104_tdata;
 wire  struct_accessed_INT_104_tvalid;
 wire  struct_accessed_INT_104_tready;

struct_access#(
.STRUCT_WIDTH(256),
.ACCESS_OFFSET(0),
.ACCESS_SIZE(32)
)struct_access_103(
	 .clk(clk), 
	 .rst(rst) ,
	//struct input
	.s_struct_axis_tdata({select_result_95_1_tdata}),
	.s_struct_axis_tvalid({select_result_95_1_tvalid}),
	.s_struct_axis_tready({select_result_95_1_tready}),
	//output val
	.m_val_axis_tdata({struct_accessed_INT_104_tdata}),
	.m_val_axis_tvalid({struct_accessed_INT_104_tvalid}),
	.m_val_axis_tready({struct_accessed_INT_104_tready})
);

//Access Struct
 wire [32-1:0] struct_accessed_INT_106_tdata;
 wire  struct_accessed_INT_106_tvalid;
 wire  struct_accessed_INT_106_tready;

struct_access#(
.STRUCT_WIDTH(256),
.ACCESS_OFFSET(128),
.ACCESS_SIZE(32)
)struct_access_105(
	 .clk(clk), 
	 .rst(rst) ,
	//struct input
	.s_struct_axis_tdata({select_result_95_2_tdata}),
	.s_struct_axis_tvalid({select_result_95_2_tvalid}),
	.s_struct_axis_tready({select_result_95_2_tready}),
	//output val
	.m_val_axis_tdata({struct_accessed_INT_106_tdata}),
	.m_val_axis_tvalid({struct_accessed_INT_106_tvalid}),
	.m_val_axis_tready({struct_accessed_INT_106_tready})
);

//Access Struct
 wire [32-1:0] struct_accessed_INT_108_tdata;
 wire  struct_accessed_INT_108_tvalid;
 wire  struct_accessed_INT_108_tready;

struct_access#(
.STRUCT_WIDTH(256),
.ACCESS_OFFSET(96),
.ACCESS_SIZE(32)
)struct_access_107(
	 .clk(clk), 
	 .rst(rst) ,
	//struct input
	.s_struct_axis_tdata({select_result_95_3_tdata}),
	.s_struct_axis_tvalid({select_result_95_3_tvalid}),
	.s_struct_axis_tready({select_result_95_3_tready}),
	//output val
	.m_val_axis_tdata({struct_accessed_INT_108_tdata}),
	.m_val_axis_tvalid({struct_accessed_INT_108_tvalid}),
	.m_val_axis_tready({struct_accessed_INT_108_tready})
);

//struct_assign_109 output struct
 wire [96-1:0] structvar_110_tdata;
 wire  structvar_110_tvalid;
 wire  structvar_110_tready;

struct_assign#(
.STRUCT_WIDTH(96),
.ASSIGN_OFFSET(0),
.ASSIGN_SIZE(32)
)struct_assign_109(
	 .clk(clk), 
	 .rst(rst) ,
	//input struct
	.s_struct_axis_tdata({inited_STRUCT_44_tdata}),
	.s_struct_axis_tvalid({inited_STRUCT_44_tvalid}),
	.s_struct_axis_tready({inited_STRUCT_44_tready}),
	//input val
	.s_assignv_axis_tdata({struct_accessed_INT_104_tdata}),
	.s_assignv_axis_tvalid({struct_accessed_INT_104_tvalid}),
	.s_assignv_axis_tready({struct_accessed_INT_104_tready}),
	//output struct
	.m_struct_axis_tdata({structvar_110_tdata}),
	.m_struct_axis_tvalid({structvar_110_tvalid}),
	.m_struct_axis_tready({structvar_110_tready})
);

//struct_assign_111 output struct
 wire [96-1:0] structvar_112_tdata;
 wire  structvar_112_tvalid;
 wire  structvar_112_tready;

struct_assign#(
.STRUCT_WIDTH(96),
.ASSIGN_OFFSET(32),
.ASSIGN_SIZE(32)
)struct_assign_111(
	 .clk(clk), 
	 .rst(rst) ,
	//input struct
	.s_struct_axis_tdata({structvar_110_tdata}),
	.s_struct_axis_tvalid({structvar_110_tvalid}),
	.s_struct_axis_tready({structvar_110_tready}),
	//input val
	.s_assignv_axis_tdata({struct_accessed_INT_106_tdata}),
	.s_assignv_axis_tvalid({struct_accessed_INT_106_tvalid}),
	.s_assignv_axis_tready({struct_accessed_INT_106_tready}),
	//output struct
	.m_struct_axis_tdata({structvar_112_tdata}),
	.m_struct_axis_tvalid({structvar_112_tvalid}),
	.m_struct_axis_tready({structvar_112_tready})
);

//struct_assign_113 output struct
 wire [96-1:0] structvar_114_tdata;
 wire  structvar_114_tvalid;
 wire  structvar_114_tready;

struct_assign#(
.STRUCT_WIDTH(96),
.ASSIGN_OFFSET(64),
.ASSIGN_SIZE(32)
)struct_assign_113(
	 .clk(clk), 
	 .rst(rst) ,
	//input struct
	.s_struct_axis_tdata({structvar_112_tdata}),
	.s_struct_axis_tvalid({structvar_112_tvalid}),
	.s_struct_axis_tready({structvar_112_tready}),
	//input val
	.s_assignv_axis_tdata({struct_accessed_INT_108_tdata}),
	.s_assignv_axis_tvalid({struct_accessed_INT_108_tvalid}),
	.s_assignv_axis_tready({struct_accessed_INT_108_tready}),
	//output struct
	.m_struct_axis_tdata({structvar_114_tdata}),
	.m_struct_axis_tvalid({structvar_114_tvalid}),
	.m_struct_axis_tready({structvar_114_tready})
);

//replicated guard condition
 wire [1-1:0] replicated_guard_cond_115_tdata;
 wire  replicated_guard_cond_115_tvalid;
 wire  replicated_guard_cond_115_tready;

//replicated guard condition
 wire [1-1:0] replicated_guard_cond_116_tdata;
 wire  replicated_guard_cond_116_tvalid;
 wire  replicated_guard_cond_116_tready;

//replicated guard condition
 wire [1-1:0] replicated_guard_cond_117_tdata;
 wire  replicated_guard_cond_117_tvalid;
 wire  replicated_guard_cond_117_tready;

//replicated guard condition
 wire [1-1:0] replicated_guard_cond_118_tdata;
 wire  replicated_guard_cond_118_tvalid;
 wire  replicated_guard_cond_118_tready;

//replicated guard condition
 wire [1-1:0] replicated_guard_cond_119_tdata;
 wire  replicated_guard_cond_119_tvalid;
 wire  replicated_guard_cond_119_tready;

guard_pred#(
.COND_WIDTH(1),
.REPLICATED_OUT_NUM(5),
.GROUND_TRUTH(1)
)guard_pred_120(
	 .clk(clk), 
	 .rst(rst) ,
	//guard condition
	.s_guard_cond_tdata({LE_65_out_INT_66_1_tdata}),
	.s_guard_cond_tvalid({LE_65_out_INT_66_1_tvalid}),
	.s_guard_cond_tready({LE_65_out_INT_66_1_tready}),
	//replicated guard condition
	.m_guard_cond_tdata({replicated_guard_cond_115_tdata,replicated_guard_cond_116_tdata,replicated_guard_cond_117_tdata,replicated_guard_cond_118_tdata,replicated_guard_cond_119_tdata}),
	.m_guard_cond_tvalid({replicated_guard_cond_115_tvalid,replicated_guard_cond_116_tvalid,replicated_guard_cond_117_tvalid,replicated_guard_cond_118_tvalid,replicated_guard_cond_119_tvalid}),
	.m_guard_cond_tready({replicated_guard_cond_115_tready,replicated_guard_cond_116_tready,replicated_guard_cond_117_tready,replicated_guard_cond_118_tready,replicated_guard_cond_119_tready})
);

//Outport Assign Src Value-- guarded
 wire [96-1:0] structvar_114_guarded_tdata;
 wire  structvar_114_guarded_tvalid;
 wire  structvar_114_guarded_tready;

guard#(
.DATA_WIDTH(96),
.IF_STREAM(0)
)guard_121(
	 .clk(clk), 
	 .rst(rst) ,
	//input val
	.s_guard_axis_tdata({structvar_114_tdata}),
	.s_guard_axis_tvalid({structvar_114_tvalid}),
	.s_guard_axis_tready({structvar_114_tready}),
	//output val
	.m_guard_axis_tdata({structvar_114_guarded_tdata}),
	.m_guard_axis_tvalid({structvar_114_guarded_tvalid}),
	.m_guard_axis_tready({structvar_114_guarded_tready}),
	//guard condition
	.s_guard_cond_tdata({replicated_guard_cond_115_tdata}),
	.s_guard_cond_tvalid({replicated_guard_cond_115_tvalid}),
	.s_guard_cond_tready({replicated_guard_cond_115_tready})
);

 assign outport_33_1_tdata = structvar_114_guarded_tdata;
 assign outport_33_1_tvalid = structvar_114_guarded_tvalid;
 assign structvar_114_guarded_tready = outport_33_1_tready;

//Outport Assign Src Value-- guarded
 wire [512-1:0] arg_29_guarded_tdata;
 wire [64-1:0] arg_29_guarded_tkeep;
 wire  arg_29_guarded_tvalid;
 wire  arg_29_guarded_tready;
 wire  arg_29_guarded_tlast;

guard#(
.DATA_WIDTH(512),
.IF_STREAM(1)
)guard_122(
	 .clk(clk), 
	 .rst(rst) ,
	//input val
	.s_guard_axis_tdata({arg_29_tdata}),
	.s_guard_axis_tkeep({arg_29_tkeep}),
	.s_guard_axis_tlast({arg_29_tlast}),
	.s_guard_axis_tvalid({arg_29_tvalid}),
	.s_guard_axis_tready({arg_29_tready}),
	//output val
	.m_guard_axis_tdata({arg_29_guarded_tdata}),
	.m_guard_axis_tkeep({arg_29_guarded_tkeep}),
	.m_guard_axis_tlast({arg_29_guarded_tlast}),
	.m_guard_axis_tvalid({arg_29_guarded_tvalid}),
	.m_guard_axis_tready({arg_29_guarded_tready}),
	//guard condition
	.s_guard_cond_tdata({replicated_guard_cond_116_tdata}),
	.s_guard_cond_tvalid({replicated_guard_cond_116_tvalid}),
	.s_guard_cond_tready({replicated_guard_cond_116_tready})
);

 assign outport_33_2_tdata = arg_29_guarded_tdata;
 assign outport_33_2_tvalid = arg_29_guarded_tvalid;
 assign arg_29_guarded_tready = outport_33_2_tready;
 assign outport_33_2_tkeep = arg_29_guarded_tkeep;
 assign outport_33_2_tlast = arg_29_guarded_tlast;

//Outport Assign Src Value-- guarded
 wire [184-1:0] arg_30_guarded_tdata;
 wire  arg_30_guarded_tvalid;
 wire  arg_30_guarded_tready;

guard#(
.DATA_WIDTH(184),
.IF_STREAM(0)
)guard_123(
	 .clk(clk), 
	 .rst(rst) ,
	//input val
	.s_guard_axis_tdata({arg_30_tdata}),
	.s_guard_axis_tvalid({arg_30_tvalid}),
	.s_guard_axis_tready({arg_30_tready}),
	//output val
	.m_guard_axis_tdata({arg_30_guarded_tdata}),
	.m_guard_axis_tvalid({arg_30_guarded_tvalid}),
	.m_guard_axis_tready({arg_30_guarded_tready}),
	//guard condition
	.s_guard_cond_tdata({replicated_guard_cond_117_tdata}),
	.s_guard_cond_tvalid({replicated_guard_cond_117_tvalid}),
	.s_guard_cond_tready({replicated_guard_cond_117_tready})
);

 assign outport_33_3_tdata = arg_30_guarded_tdata;
 assign outport_33_3_tvalid = arg_30_guarded_tvalid;
 assign arg_30_guarded_tready = outport_33_3_tready;

//Outport Assign Src Value-- guarded
 wire [112-1:0] arg_31_guarded_tdata;
 wire  arg_31_guarded_tvalid;
 wire  arg_31_guarded_tready;

guard#(
.DATA_WIDTH(112),
.IF_STREAM(0)
)guard_124(
	 .clk(clk), 
	 .rst(rst) ,
	//input val
	.s_guard_axis_tdata({arg_31_tdata}),
	.s_guard_axis_tvalid({arg_31_tvalid}),
	.s_guard_axis_tready({arg_31_tready}),
	//output val
	.m_guard_axis_tdata({arg_31_guarded_tdata}),
	.m_guard_axis_tvalid({arg_31_guarded_tvalid}),
	.m_guard_axis_tready({arg_31_guarded_tready}),
	//guard condition
	.s_guard_cond_tdata({replicated_guard_cond_118_tdata}),
	.s_guard_cond_tvalid({replicated_guard_cond_118_tvalid}),
	.s_guard_cond_tready({replicated_guard_cond_118_tready})
);

 assign outport_33_4_tdata = arg_31_guarded_tdata;
 assign outport_33_4_tvalid = arg_31_guarded_tvalid;
 assign arg_31_guarded_tready = outport_33_4_tready;

//Outport Assign Src Value-- guarded
 wire [160-1:0] arg_32_guarded_tdata;
 wire  arg_32_guarded_tvalid;
 wire  arg_32_guarded_tready;

guard#(
.DATA_WIDTH(160),
.IF_STREAM(0)
)guard_125(
	 .clk(clk), 
	 .rst(rst) ,
	//input val
	.s_guard_axis_tdata({arg_32_tdata}),
	.s_guard_axis_tvalid({arg_32_tvalid}),
	.s_guard_axis_tready({arg_32_tready}),
	//output val
	.m_guard_axis_tdata({arg_32_guarded_tdata}),
	.m_guard_axis_tvalid({arg_32_guarded_tvalid}),
	.m_guard_axis_tready({arg_32_guarded_tready}),
	//guard condition
	.s_guard_cond_tdata({replicated_guard_cond_119_tdata}),
	.s_guard_cond_tvalid({replicated_guard_cond_119_tvalid}),
	.s_guard_cond_tready({replicated_guard_cond_119_tready})
);

 assign outport_33_5_tdata = arg_32_guarded_tdata;
 assign outport_33_5_tvalid = arg_32_guarded_tvalid;
 assign arg_32_guarded_tready = outport_33_5_tready;


endmodule
