module __handler_NET_SEND#()
(
	 input  wire clk, 
	 input  wire rst,
	//input ports BUF
	input wire [512-1:0] arg1_tdata ,
	input wire [64-1:0] arg1_tkeep ,
	input wire  arg1_tlast ,
	input wire  arg1_tvalid ,
	output wire  arg1_tready
);

endmodule
